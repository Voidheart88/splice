Vin 1 0 10
R1 1 2 1000
R2 2 0 1000
E1 3 0 2 0 2.0
G1 3 4 2 0 0.01
.op
.end