*Test*
.model diode D()
V1 N0 0 10
R1 N0 N1 10
D1 N1 0 diode
R2 N1 N2 10
D2 N2 0 diode
R3 N2 N3 10
D3 N3 0 diode
R4 N3 N4 10
D4 N4 0 diode
R5 N4 N5 10
D5 N5 0 diode
R6 N5 N6 10
D6 N6 0 diode
R7 N6 N7 10
D7 N7 0 diode
R8 N7 N8 10
D8 N8 0 diode
R9 N8 N9 10
D9 N9 0 diode
R10 N9 N10 10
D10 N10 0 diode
R11 N10 N11 10
D11 N11 0 diode
R12 N11 N12 10
D12 N12 0 diode
R13 N12 N13 10
D13 N13 0 diode
R14 N13 N14 10
D14 N14 0 diode
R15 N14 N15 10
D15 N15 0 diode
R16 N15 N16 10
D16 N16 0 diode
R17 N16 N17 10
D17 N17 0 diode
R18 N17 N18 10
D18 N18 0 diode
R19 N18 N19 10
D19 N19 0 diode
R20 N19 N20 10
D20 N20 0 diode
R21 N20 N21 10
D21 N21 0 diode
R22 N21 N22 10
D22 N22 0 diode
R23 N22 N23 10
D23 N23 0 diode
R24 N23 N24 10
D24 N24 0 diode
R25 N24 N25 10
D25 N25 0 diode
R26 N25 N26 10
D26 N26 0 diode
R27 N26 N27 10
D27 N27 0 diode
R28 N27 N28 10
D28 N28 0 diode
R29 N28 N29 10
D29 N29 0 diode
R30 N29 N30 10
D30 N30 0 diode
R31 N30 N31 10
D31 N31 0 diode
R32 N31 N32 10
D32 N32 0 diode
R33 N32 N33 10
D33 N33 0 diode
R34 N33 N34 10
D34 N34 0 diode
R35 N34 N35 10
D35 N35 0 diode
R36 N35 N36 10
D36 N36 0 diode
R37 N36 N37 10
D37 N37 0 diode
R38 N37 N38 10
D38 N38 0 diode
R39 N38 N39 10
D39 N39 0 diode
R40 N39 N40 10
D40 N40 0 diode
R41 N40 N41 10
D41 N41 0 diode
R42 N41 N42 10
D42 N42 0 diode
R43 N42 N43 10
D43 N43 0 diode
R44 N43 N44 10
D44 N44 0 diode
R45 N44 N45 10
D45 N45 0 diode
R46 N45 N46 10
D46 N46 0 diode
R47 N46 N47 10
D47 N47 0 diode
R48 N47 N48 10
D48 N48 0 diode
R49 N48 N49 10
D49 N49 0 diode
R50 N49 N50 10
D50 N50 0 diode
R51 N50 N51 10
D51 N51 0 diode
R52 N51 N52 10
D52 N52 0 diode
R53 N52 N53 10
D53 N53 0 diode
R54 N53 N54 10
D54 N54 0 diode
R55 N54 N55 10
D55 N55 0 diode
R56 N55 N56 10
D56 N56 0 diode
R57 N56 N57 10
D57 N57 0 diode
R58 N57 N58 10
D58 N58 0 diode
R59 N58 N59 10
D59 N59 0 diode
R60 N59 N60 10
D60 N60 0 diode
R61 N60 N61 10
D61 N61 0 diode
R62 N61 N62 10
D62 N62 0 diode
R63 N62 N63 10
D63 N63 0 diode
R64 N63 N64 10
D64 N64 0 diode
R65 N64 N65 10
D65 N65 0 diode
R66 N65 N66 10
D66 N66 0 diode
R67 N66 N67 10
D67 N67 0 diode
R68 N67 N68 10
D68 N68 0 diode
R69 N68 N69 10
D69 N69 0 diode
R70 N69 N70 10
D70 N70 0 diode
R71 N70 N71 10
D71 N71 0 diode
R72 N71 N72 10
D72 N72 0 diode
R73 N72 N73 10
D73 N73 0 diode
R74 N73 N74 10
D74 N74 0 diode
R75 N74 N75 10
D75 N75 0 diode
R76 N75 N76 10
D76 N76 0 diode
R77 N76 N77 10
D77 N77 0 diode
R78 N77 N78 10
D78 N78 0 diode
R79 N78 N79 10
D79 N79 0 diode
R80 N79 N80 10
D80 N80 0 diode
R81 N80 N81 10
D81 N81 0 diode
R82 N81 N82 10
D82 N82 0 diode
R83 N82 N83 10
D83 N83 0 diode
R84 N83 N84 10
D84 N84 0 diode
R85 N84 N85 10
D85 N85 0 diode
R86 N85 N86 10
D86 N86 0 diode
R87 N86 N87 10
D87 N87 0 diode
R88 N87 N88 10
D88 N88 0 diode
R89 N88 N89 10
D89 N89 0 diode
R90 N89 N90 10
D90 N90 0 diode
R91 N90 N91 10
D91 N91 0 diode
R92 N91 N92 10
D92 N92 0 diode
R93 N92 N93 10
D93 N93 0 diode
R94 N93 N94 10
D94 N94 0 diode
R95 N94 N95 10
D95 N95 0 diode
R96 N95 N96 10
D96 N96 0 diode
R97 N96 N97 10
D97 N97 0 diode
R98 N97 N98 10
D98 N98 0 diode
R99 N98 N99 10
D99 N99 0 diode
R100 N99 N100 10
D100 N100 0 diode
R101 N100 N101 10
D101 N101 0 diode
R102 N101 N102 10
D102 N102 0 diode
R103 N102 N103 10
D103 N103 0 diode
R104 N103 N104 10
D104 N104 0 diode
R105 N104 N105 10
D105 N105 0 diode
R106 N105 N106 10
D106 N106 0 diode
R107 N106 N107 10
D107 N107 0 diode
R108 N107 N108 10
D108 N108 0 diode
R109 N108 N109 10
D109 N109 0 diode
R110 N109 N110 10
D110 N110 0 diode
R111 N110 N111 10
D111 N111 0 diode
R112 N111 N112 10
D112 N112 0 diode
R113 N112 N113 10
D113 N113 0 diode
R114 N113 N114 10
D114 N114 0 diode
R115 N114 N115 10
D115 N115 0 diode
R116 N115 N116 10
D116 N116 0 diode
R117 N116 N117 10
D117 N117 0 diode
R118 N117 N118 10
D118 N118 0 diode
R119 N118 N119 10
D119 N119 0 diode
R120 N119 N120 10
D120 N120 0 diode
R121 N120 N121 10
D121 N121 0 diode
R122 N121 N122 10
D122 N122 0 diode
R123 N122 N123 10
D123 N123 0 diode
R124 N123 N124 10
D124 N124 0 diode
R125 N124 N125 10
D125 N125 0 diode
R126 N125 N126 10
D126 N126 0 diode
R127 N126 N127 10
D127 N127 0 diode
R128 N127 N128 10
D128 N128 0 diode
R129 N128 N129 10
D129 N129 0 diode
R130 N129 N130 10
D130 N130 0 diode
R131 N130 N131 10
D131 N131 0 diode
R132 N131 N132 10
D132 N132 0 diode
R133 N132 N133 10
D133 N133 0 diode
R134 N133 N134 10
D134 N134 0 diode
R135 N134 N135 10
D135 N135 0 diode
R136 N135 N136 10
D136 N136 0 diode
R137 N136 N137 10
D137 N137 0 diode
R138 N137 N138 10
D138 N138 0 diode
R139 N138 N139 10
D139 N139 0 diode
R140 N139 N140 10
D140 N140 0 diode
R141 N140 N141 10
D141 N141 0 diode
R142 N141 N142 10
D142 N142 0 diode
R143 N142 N143 10
D143 N143 0 diode
R144 N143 N144 10
D144 N144 0 diode
R145 N144 N145 10
D145 N145 0 diode
R146 N145 N146 10
D146 N146 0 diode
R147 N146 N147 10
D147 N147 0 diode
R148 N147 N148 10
D148 N148 0 diode
R149 N148 N149 10
D149 N149 0 diode
R150 N149 N150 10
D150 N150 0 diode
R151 N150 N151 10
D151 N151 0 diode
R152 N151 N152 10
D152 N152 0 diode
R153 N152 N153 10
D153 N153 0 diode
R154 N153 N154 10
D154 N154 0 diode
R155 N154 N155 10
D155 N155 0 diode
R156 N155 N156 10
D156 N156 0 diode
R157 N156 N157 10
D157 N157 0 diode
R158 N157 N158 10
D158 N158 0 diode
R159 N158 N159 10
D159 N159 0 diode
R160 N159 N160 10
D160 N160 0 diode
R161 N160 N161 10
D161 N161 0 diode
R162 N161 N162 10
D162 N162 0 diode
R163 N162 N163 10
D163 N163 0 diode
R164 N163 N164 10
D164 N164 0 diode
R165 N164 N165 10
D165 N165 0 diode
R166 N165 N166 10
D166 N166 0 diode
R167 N166 N167 10
D167 N167 0 diode
R168 N167 N168 10
D168 N168 0 diode
R169 N168 N169 10
D169 N169 0 diode
R170 N169 N170 10
D170 N170 0 diode
R171 N170 N171 10
D171 N171 0 diode
R172 N171 N172 10
D172 N172 0 diode
R173 N172 N173 10
D173 N173 0 diode
R174 N173 N174 10
D174 N174 0 diode
R175 N174 N175 10
D175 N175 0 diode
R176 N175 N176 10
D176 N176 0 diode
R177 N176 N177 10
D177 N177 0 diode
R178 N177 N178 10
D178 N178 0 diode
R179 N178 N179 10
D179 N179 0 diode
R180 N179 N180 10
D180 N180 0 diode
R181 N180 N181 10
D181 N181 0 diode
R182 N181 N182 10
D182 N182 0 diode
R183 N182 N183 10
D183 N183 0 diode
R184 N183 N184 10
D184 N184 0 diode
R185 N184 N185 10
D185 N185 0 diode
R186 N185 N186 10
D186 N186 0 diode
R187 N186 N187 10
D187 N187 0 diode
R188 N187 N188 10
D188 N188 0 diode
R189 N188 N189 10
D189 N189 0 diode
R190 N189 N190 10
D190 N190 0 diode
R191 N190 N191 10
D191 N191 0 diode
R192 N191 N192 10
D192 N192 0 diode
R193 N192 N193 10
D193 N193 0 diode
R194 N193 N194 10
D194 N194 0 diode
R195 N194 N195 10
D195 N195 0 diode
R196 N195 N196 10
D196 N196 0 diode
R197 N196 N197 10
D197 N197 0 diode
R198 N197 N198 10
D198 N198 0 diode
R199 N198 N199 10
D199 N199 0 diode
R200 N199 N200 10
D200 N200 0 diode
R201 N200 N201 10
D201 N201 0 diode
R202 N201 N202 10
D202 N202 0 diode
R203 N202 N203 10
D203 N203 0 diode
R204 N203 N204 10
D204 N204 0 diode
R205 N204 N205 10
D205 N205 0 diode
R206 N205 N206 10
D206 N206 0 diode
R207 N206 N207 10
D207 N207 0 diode
R208 N207 N208 10
D208 N208 0 diode
R209 N208 N209 10
D209 N209 0 diode
R210 N209 N210 10
D210 N210 0 diode
R211 N210 N211 10
D211 N211 0 diode
R212 N211 N212 10
D212 N212 0 diode
R213 N212 N213 10
D213 N213 0 diode
R214 N213 N214 10
D214 N214 0 diode
R215 N214 N215 10
D215 N215 0 diode
R216 N215 N216 10
D216 N216 0 diode
R217 N216 N217 10
D217 N217 0 diode
R218 N217 N218 10
D218 N218 0 diode
R219 N218 N219 10
D219 N219 0 diode
R220 N219 N220 10
D220 N220 0 diode
R221 N220 N221 10
D221 N221 0 diode
R222 N221 N222 10
D222 N222 0 diode
R223 N222 N223 10
D223 N223 0 diode
R224 N223 N224 10
D224 N224 0 diode
R225 N224 N225 10
D225 N225 0 diode
R226 N225 N226 10
D226 N226 0 diode
R227 N226 N227 10
D227 N227 0 diode
R228 N227 N228 10
D228 N228 0 diode
R229 N228 N229 10
D229 N229 0 diode
R230 N229 N230 10
D230 N230 0 diode
R231 N230 N231 10
D231 N231 0 diode
R232 N231 N232 10
D232 N232 0 diode
R233 N232 N233 10
D233 N233 0 diode
R234 N233 N234 10
D234 N234 0 diode
R235 N234 N235 10
D235 N235 0 diode
R236 N235 N236 10
D236 N236 0 diode
R237 N236 N237 10
D237 N237 0 diode
R238 N237 N238 10
D238 N238 0 diode
R239 N238 N239 10
D239 N239 0 diode
R240 N239 N240 10
D240 N240 0 diode
R241 N240 N241 10
D241 N241 0 diode
R242 N241 N242 10
D242 N242 0 diode
R243 N242 N243 10
D243 N243 0 diode
R244 N243 N244 10
D244 N244 0 diode
R245 N244 N245 10
D245 N245 0 diode
R246 N245 N246 10
D246 N246 0 diode
R247 N246 N247 10
D247 N247 0 diode
R248 N247 N248 10
D248 N248 0 diode
R249 N248 N249 10
D249 N249 0 diode
R250 N249 N250 10
D250 N250 0 diode
R251 N250 N251 10
D251 N251 0 diode
R252 N251 N252 10
D252 N252 0 diode
R253 N252 N253 10
D253 N253 0 diode
R254 N253 N254 10
D254 N254 0 diode
R255 N254 N255 10
D255 N255 0 diode
R256 N255 N256 10
D256 N256 0 diode
R257 N256 N257 10
D257 N257 0 diode
R258 N257 N258 10
D258 N258 0 diode
R259 N258 N259 10
D259 N259 0 diode
R260 N259 N260 10
D260 N260 0 diode
R261 N260 N261 10
D261 N261 0 diode
R262 N261 N262 10
D262 N262 0 diode
R263 N262 N263 10
D263 N263 0 diode
R264 N263 N264 10
D264 N264 0 diode
R265 N264 N265 10
D265 N265 0 diode
R266 N265 N266 10
D266 N266 0 diode
R267 N266 N267 10
D267 N267 0 diode
R268 N267 N268 10
D268 N268 0 diode
R269 N268 N269 10
D269 N269 0 diode
R270 N269 N270 10
D270 N270 0 diode
R271 N270 N271 10
D271 N271 0 diode
R272 N271 N272 10
D272 N272 0 diode
R273 N272 N273 10
D273 N273 0 diode
R274 N273 N274 10
D274 N274 0 diode
R275 N274 N275 10
D275 N275 0 diode
R276 N275 N276 10
D276 N276 0 diode
R277 N276 N277 10
D277 N277 0 diode
R278 N277 N278 10
D278 N278 0 diode
R279 N278 N279 10
D279 N279 0 diode
R280 N279 N280 10
D280 N280 0 diode
R281 N280 N281 10
D281 N281 0 diode
R282 N281 N282 10
D282 N282 0 diode
R283 N282 N283 10
D283 N283 0 diode
R284 N283 N284 10
D284 N284 0 diode
R285 N284 N285 10
D285 N285 0 diode
R286 N285 N286 10
D286 N286 0 diode
R287 N286 N287 10
D287 N287 0 diode
R288 N287 N288 10
D288 N288 0 diode
R289 N288 N289 10
D289 N289 0 diode
R290 N289 N290 10
D290 N290 0 diode
R291 N290 N291 10
D291 N291 0 diode
R292 N291 N292 10
D292 N292 0 diode
R293 N292 N293 10
D293 N293 0 diode
R294 N293 N294 10
D294 N294 0 diode
R295 N294 N295 10
D295 N295 0 diode
R296 N295 N296 10
D296 N296 0 diode
R297 N296 N297 10
D297 N297 0 diode
R298 N297 N298 10
D298 N298 0 diode
R299 N298 N299 10
D299 N299 0 diode
R300 N299 N300 10
D300 N300 0 diode
R301 N300 N301 10
D301 N301 0 diode
R302 N301 N302 10
D302 N302 0 diode
R303 N302 N303 10
D303 N303 0 diode
R304 N303 N304 10
D304 N304 0 diode
R305 N304 N305 10
D305 N305 0 diode
R306 N305 N306 10
D306 N306 0 diode
R307 N306 N307 10
D307 N307 0 diode
R308 N307 N308 10
D308 N308 0 diode
R309 N308 N309 10
D309 N309 0 diode
R310 N309 N310 10
D310 N310 0 diode
R311 N310 N311 10
D311 N311 0 diode
R312 N311 N312 10
D312 N312 0 diode
R313 N312 N313 10
D313 N313 0 diode
R314 N313 N314 10
D314 N314 0 diode
R315 N314 N315 10
D315 N315 0 diode
R316 N315 N316 10
D316 N316 0 diode
R317 N316 N317 10
D317 N317 0 diode
R318 N317 N318 10
D318 N318 0 diode
R319 N318 N319 10
D319 N319 0 diode
R320 N319 N320 10
D320 N320 0 diode
R321 N320 N321 10
D321 N321 0 diode
R322 N321 N322 10
D322 N322 0 diode
R323 N322 N323 10
D323 N323 0 diode
R324 N323 N324 10
D324 N324 0 diode
R325 N324 N325 10
D325 N325 0 diode
R326 N325 N326 10
D326 N326 0 diode
R327 N326 N327 10
D327 N327 0 diode
R328 N327 N328 10
D328 N328 0 diode
R329 N328 N329 10
D329 N329 0 diode
R330 N329 N330 10
D330 N330 0 diode
R331 N330 N331 10
D331 N331 0 diode
R332 N331 N332 10
D332 N332 0 diode
R333 N332 N333 10
D333 N333 0 diode
R334 N333 N334 10
D334 N334 0 diode
R335 N334 N335 10
D335 N335 0 diode
R336 N335 N336 10
D336 N336 0 diode
R337 N336 N337 10
D337 N337 0 diode
R338 N337 N338 10
D338 N338 0 diode
R339 N338 N339 10
D339 N339 0 diode
R340 N339 N340 10
D340 N340 0 diode
R341 N340 N341 10
D341 N341 0 diode
R342 N341 N342 10
D342 N342 0 diode
R343 N342 N343 10
D343 N343 0 diode
R344 N343 N344 10
D344 N344 0 diode
R345 N344 N345 10
D345 N345 0 diode
R346 N345 N346 10
D346 N346 0 diode
R347 N346 N347 10
D347 N347 0 diode
R348 N347 N348 10
D348 N348 0 diode
R349 N348 N349 10
D349 N349 0 diode
R350 N349 N350 10
D350 N350 0 diode
R351 N350 N351 10
D351 N351 0 diode
R352 N351 N352 10
D352 N352 0 diode
R353 N352 N353 10
D353 N353 0 diode
R354 N353 N354 10
D354 N354 0 diode
R355 N354 N355 10
D355 N355 0 diode
R356 N355 N356 10
D356 N356 0 diode
R357 N356 N357 10
D357 N357 0 diode
R358 N357 N358 10
D358 N358 0 diode
R359 N358 N359 10
D359 N359 0 diode
R360 N359 N360 10
D360 N360 0 diode
R361 N360 N361 10
D361 N361 0 diode
R362 N361 N362 10
D362 N362 0 diode
R363 N362 N363 10
D363 N363 0 diode
R364 N363 N364 10
D364 N364 0 diode
R365 N364 N365 10
D365 N365 0 diode
R366 N365 N366 10
D366 N366 0 diode
R367 N366 N367 10
D367 N367 0 diode
R368 N367 N368 10
D368 N368 0 diode
R369 N368 N369 10
D369 N369 0 diode
R370 N369 N370 10
D370 N370 0 diode
R371 N370 N371 10
D371 N371 0 diode
R372 N371 N372 10
D372 N372 0 diode
R373 N372 N373 10
D373 N373 0 diode
R374 N373 N374 10
D374 N374 0 diode
R375 N374 N375 10
D375 N375 0 diode
R376 N375 N376 10
D376 N376 0 diode
R377 N376 N377 10
D377 N377 0 diode
R378 N377 N378 10
D378 N378 0 diode
R379 N378 N379 10
D379 N379 0 diode
R380 N379 N380 10
D380 N380 0 diode
R381 N380 N381 10
D381 N381 0 diode
R382 N381 N382 10
D382 N382 0 diode
R383 N382 N383 10
D383 N383 0 diode
R384 N383 N384 10
D384 N384 0 diode
R385 N384 N385 10
D385 N385 0 diode
R386 N385 N386 10
D386 N386 0 diode
R387 N386 N387 10
D387 N387 0 diode
R388 N387 N388 10
D388 N388 0 diode
R389 N388 N389 10
D389 N389 0 diode
R390 N389 N390 10
D390 N390 0 diode
R391 N390 N391 10
D391 N391 0 diode
R392 N391 N392 10
D392 N392 0 diode
R393 N392 N393 10
D393 N393 0 diode
R394 N393 N394 10
D394 N394 0 diode
R395 N394 N395 10
D395 N395 0 diode
R396 N395 N396 10
D396 N396 0 diode
R397 N396 N397 10
D397 N397 0 diode
R398 N397 N398 10
D398 N398 0 diode
R399 N398 N399 10
D399 N399 0 diode
R400 N399 N400 10
D400 N400 0 diode
R401 N400 N401 10
D401 N401 0 diode
R402 N401 N402 10
D402 N402 0 diode
R403 N402 N403 10
D403 N403 0 diode
R404 N403 N404 10
D404 N404 0 diode
R405 N404 N405 10
D405 N405 0 diode
R406 N405 N406 10
D406 N406 0 diode
R407 N406 N407 10
D407 N407 0 diode
R408 N407 N408 10
D408 N408 0 diode
R409 N408 N409 10
D409 N409 0 diode
R410 N409 N410 10
D410 N410 0 diode
R411 N410 N411 10
D411 N411 0 diode
R412 N411 N412 10
D412 N412 0 diode
R413 N412 N413 10
D413 N413 0 diode
R414 N413 N414 10
D414 N414 0 diode
R415 N414 N415 10
D415 N415 0 diode
R416 N415 N416 10
D416 N416 0 diode
R417 N416 N417 10
D417 N417 0 diode
R418 N417 N418 10
D418 N418 0 diode
R419 N418 N419 10
D419 N419 0 diode
R420 N419 N420 10
D420 N420 0 diode
R421 N420 N421 10
D421 N421 0 diode
R422 N421 N422 10
D422 N422 0 diode
R423 N422 N423 10
D423 N423 0 diode
R424 N423 N424 10
D424 N424 0 diode
R425 N424 N425 10
D425 N425 0 diode
R426 N425 N426 10
D426 N426 0 diode
R427 N426 N427 10
D427 N427 0 diode
R428 N427 N428 10
D428 N428 0 diode
R429 N428 N429 10
D429 N429 0 diode
R430 N429 N430 10
D430 N430 0 diode
R431 N430 N431 10
D431 N431 0 diode
R432 N431 N432 10
D432 N432 0 diode
R433 N432 N433 10
D433 N433 0 diode
R434 N433 N434 10
D434 N434 0 diode
R435 N434 N435 10
D435 N435 0 diode
R436 N435 N436 10
D436 N436 0 diode
R437 N436 N437 10
D437 N437 0 diode
R438 N437 N438 10
D438 N438 0 diode
R439 N438 N439 10
D439 N439 0 diode
R440 N439 N440 10
D440 N440 0 diode
R441 N440 N441 10
D441 N441 0 diode
R442 N441 N442 10
D442 N442 0 diode
R443 N442 N443 10
D443 N443 0 diode
R444 N443 N444 10
D444 N444 0 diode
R445 N444 N445 10
D445 N445 0 diode
R446 N445 N446 10
D446 N446 0 diode
R447 N446 N447 10
D447 N447 0 diode
R448 N447 N448 10
D448 N448 0 diode
R449 N448 N449 10
D449 N449 0 diode
R450 N449 N450 10
D450 N450 0 diode
R451 N450 N451 10
D451 N451 0 diode
R452 N451 N452 10
D452 N452 0 diode
R453 N452 N453 10
D453 N453 0 diode
R454 N453 N454 10
D454 N454 0 diode
R455 N454 N455 10
D455 N455 0 diode
R456 N455 N456 10
D456 N456 0 diode
R457 N456 N457 10
D457 N457 0 diode
R458 N457 N458 10
D458 N458 0 diode
R459 N458 N459 10
D459 N459 0 diode
R460 N459 N460 10
D460 N460 0 diode
R461 N460 N461 10
D461 N461 0 diode
R462 N461 N462 10
D462 N462 0 diode
R463 N462 N463 10
D463 N463 0 diode
R464 N463 N464 10
D464 N464 0 diode
R465 N464 N465 10
D465 N465 0 diode
R466 N465 N466 10
D466 N466 0 diode
R467 N466 N467 10
D467 N467 0 diode
R468 N467 N468 10
D468 N468 0 diode
R469 N468 N469 10
D469 N469 0 diode
R470 N469 N470 10
D470 N470 0 diode
R471 N470 N471 10
D471 N471 0 diode
R472 N471 N472 10
D472 N472 0 diode
R473 N472 N473 10
D473 N473 0 diode
R474 N473 N474 10
D474 N474 0 diode
R475 N474 N475 10
D475 N475 0 diode
R476 N475 N476 10
D476 N476 0 diode
R477 N476 N477 10
D477 N477 0 diode
R478 N477 N478 10
D478 N478 0 diode
R479 N478 N479 10
D479 N479 0 diode
R480 N479 N480 10
D480 N480 0 diode
R481 N480 N481 10
D481 N481 0 diode
R482 N481 N482 10
D482 N482 0 diode
R483 N482 N483 10
D483 N483 0 diode
R484 N483 N484 10
D484 N484 0 diode
R485 N484 N485 10
D485 N485 0 diode
R486 N485 N486 10
D486 N486 0 diode
R487 N486 N487 10
D487 N487 0 diode
R488 N487 N488 10
D488 N488 0 diode
R489 N488 N489 10
D489 N489 0 diode
R490 N489 N490 10
D490 N490 0 diode
R491 N490 N491 10
D491 N491 0 diode
R492 N491 N492 10
D492 N492 0 diode
R493 N492 N493 10
D493 N493 0 diode
R494 N493 N494 10
D494 N494 0 diode
R495 N494 N495 10
D495 N495 0 diode
R496 N495 N496 10
D496 N496 0 diode
R497 N496 N497 10
D497 N497 0 diode
R498 N497 N498 10
D498 N498 0 diode
R499 N498 N499 10
D499 N499 0 diode
R500 N499 N500 10
D500 N500 0 diode
R501 N500 N501 10
D501 N501 0 diode
R502 N501 N502 10
D502 N502 0 diode
R503 N502 N503 10
D503 N503 0 diode
R504 N503 N504 10
D504 N504 0 diode
R505 N504 N505 10
D505 N505 0 diode
R506 N505 N506 10
D506 N506 0 diode
R507 N506 N507 10
D507 N507 0 diode
R508 N507 N508 10
D508 N508 0 diode
R509 N508 N509 10
D509 N509 0 diode
R510 N509 N510 10
D510 N510 0 diode
R511 N510 N511 10
D511 N511 0 diode
R512 N511 N512 10
D512 N512 0 diode
R513 N512 N513 10
D513 N513 0 diode
R514 N513 N514 10
D514 N514 0 diode
R515 N514 N515 10
D515 N515 0 diode
R516 N515 N516 10
D516 N516 0 diode
R517 N516 N517 10
D517 N517 0 diode
R518 N517 N518 10
D518 N518 0 diode
R519 N518 N519 10
D519 N519 0 diode
R520 N519 N520 10
D520 N520 0 diode
R521 N520 N521 10
D521 N521 0 diode
R522 N521 N522 10
D522 N522 0 diode
R523 N522 N523 10
D523 N523 0 diode
R524 N523 N524 10
D524 N524 0 diode
R525 N524 N525 10
D525 N525 0 diode
R526 N525 N526 10
D526 N526 0 diode
R527 N526 N527 10
D527 N527 0 diode
R528 N527 N528 10
D528 N528 0 diode
R529 N528 N529 10
D529 N529 0 diode
R530 N529 N530 10
D530 N530 0 diode
R531 N530 N531 10
D531 N531 0 diode
R532 N531 N532 10
D532 N532 0 diode
R533 N532 N533 10
D533 N533 0 diode
R534 N533 N534 10
D534 N534 0 diode
R535 N534 N535 10
D535 N535 0 diode
R536 N535 N536 10
D536 N536 0 diode
R537 N536 N537 10
D537 N537 0 diode
R538 N537 N538 10
D538 N538 0 diode
R539 N538 N539 10
D539 N539 0 diode
R540 N539 N540 10
D540 N540 0 diode
R541 N540 N541 10
D541 N541 0 diode
R542 N541 N542 10
D542 N542 0 diode
R543 N542 N543 10
D543 N543 0 diode
R544 N543 N544 10
D544 N544 0 diode
R545 N544 N545 10
D545 N545 0 diode
R546 N545 N546 10
D546 N546 0 diode
R547 N546 N547 10
D547 N547 0 diode
R548 N547 N548 10
D548 N548 0 diode
R549 N548 N549 10
D549 N549 0 diode
R550 N549 N550 10
D550 N550 0 diode
R551 N550 N551 10
D551 N551 0 diode
R552 N551 N552 10
D552 N552 0 diode
R553 N552 N553 10
D553 N553 0 diode
R554 N553 N554 10
D554 N554 0 diode
R555 N554 N555 10
D555 N555 0 diode
R556 N555 N556 10
D556 N556 0 diode
R557 N556 N557 10
D557 N557 0 diode
R558 N557 N558 10
D558 N558 0 diode
R559 N558 N559 10
D559 N559 0 diode
R560 N559 N560 10
D560 N560 0 diode
R561 N560 N561 10
D561 N561 0 diode
R562 N561 N562 10
D562 N562 0 diode
R563 N562 N563 10
D563 N563 0 diode
R564 N563 N564 10
D564 N564 0 diode
R565 N564 N565 10
D565 N565 0 diode
R566 N565 N566 10
D566 N566 0 diode
R567 N566 N567 10
D567 N567 0 diode
R568 N567 N568 10
D568 N568 0 diode
R569 N568 N569 10
D569 N569 0 diode
R570 N569 N570 10
D570 N570 0 diode
R571 N570 N571 10
D571 N571 0 diode
R572 N571 N572 10
D572 N572 0 diode
R573 N572 N573 10
D573 N573 0 diode
R574 N573 N574 10
D574 N574 0 diode
R575 N574 N575 10
D575 N575 0 diode
R576 N575 N576 10
D576 N576 0 diode
R577 N576 N577 10
D577 N577 0 diode
R578 N577 N578 10
D578 N578 0 diode
R579 N578 N579 10
D579 N579 0 diode
R580 N579 N580 10
D580 N580 0 diode
R581 N580 N581 10
D581 N581 0 diode
R582 N581 N582 10
D582 N582 0 diode
R583 N582 N583 10
D583 N583 0 diode
R584 N583 N584 10
D584 N584 0 diode
R585 N584 N585 10
D585 N585 0 diode
R586 N585 N586 10
D586 N586 0 diode
R587 N586 N587 10
D587 N587 0 diode
R588 N587 N588 10
D588 N588 0 diode
R589 N588 N589 10
D589 N589 0 diode
R590 N589 N590 10
D590 N590 0 diode
R591 N590 N591 10
D591 N591 0 diode
R592 N591 N592 10
D592 N592 0 diode
R593 N592 N593 10
D593 N593 0 diode
R594 N593 N594 10
D594 N594 0 diode
R595 N594 N595 10
D595 N595 0 diode
R596 N595 N596 10
D596 N596 0 diode
R597 N596 N597 10
D597 N597 0 diode
R598 N597 N598 10
D598 N598 0 diode
R599 N598 N599 10
D599 N599 0 diode
R600 N599 N600 10
D600 N600 0 diode
R601 N600 N601 10
D601 N601 0 diode
R602 N601 N602 10
D602 N602 0 diode
R603 N602 N603 10
D603 N603 0 diode
R604 N603 N604 10
D604 N604 0 diode
R605 N604 N605 10
D605 N605 0 diode
R606 N605 N606 10
D606 N606 0 diode
R607 N606 N607 10
D607 N607 0 diode
R608 N607 N608 10
D608 N608 0 diode
R609 N608 N609 10
D609 N609 0 diode
R610 N609 N610 10
D610 N610 0 diode
R611 N610 N611 10
D611 N611 0 diode
R612 N611 N612 10
D612 N612 0 diode
R613 N612 N613 10
D613 N613 0 diode
R614 N613 N614 10
D614 N614 0 diode
R615 N614 N615 10
D615 N615 0 diode
R616 N615 N616 10
D616 N616 0 diode
R617 N616 N617 10
D617 N617 0 diode
R618 N617 N618 10
D618 N618 0 diode
R619 N618 N619 10
D619 N619 0 diode
R620 N619 N620 10
D620 N620 0 diode
R621 N620 N621 10
D621 N621 0 diode
R622 N621 N622 10
D622 N622 0 diode
R623 N622 N623 10
D623 N623 0 diode
R624 N623 N624 10
D624 N624 0 diode
R625 N624 N625 10
D625 N625 0 diode
R626 N625 N626 10
D626 N626 0 diode
R627 N626 N627 10
D627 N627 0 diode
R628 N627 N628 10
D628 N628 0 diode
R629 N628 N629 10
D629 N629 0 diode
R630 N629 N630 10
D630 N630 0 diode
R631 N630 N631 10
D631 N631 0 diode
R632 N631 N632 10
D632 N632 0 diode
R633 N632 N633 10
D633 N633 0 diode
R634 N633 N634 10
D634 N634 0 diode
R635 N634 N635 10
D635 N635 0 diode
R636 N635 N636 10
D636 N636 0 diode
R637 N636 N637 10
D637 N637 0 diode
R638 N637 N638 10
D638 N638 0 diode
R639 N638 N639 10
D639 N639 0 diode
R640 N639 N640 10
D640 N640 0 diode
R641 N640 N641 10
D641 N641 0 diode
R642 N641 N642 10
D642 N642 0 diode
R643 N642 N643 10
D643 N643 0 diode
R644 N643 N644 10
D644 N644 0 diode
R645 N644 N645 10
D645 N645 0 diode
R646 N645 N646 10
D646 N646 0 diode
R647 N646 N647 10
D647 N647 0 diode
R648 N647 N648 10
D648 N648 0 diode
R649 N648 N649 10
D649 N649 0 diode
R650 N649 N650 10
D650 N650 0 diode
R651 N650 N651 10
D651 N651 0 diode
R652 N651 N652 10
D652 N652 0 diode
R653 N652 N653 10
D653 N653 0 diode
R654 N653 N654 10
D654 N654 0 diode
R655 N654 N655 10
D655 N655 0 diode
R656 N655 N656 10
D656 N656 0 diode
R657 N656 N657 10
D657 N657 0 diode
R658 N657 N658 10
D658 N658 0 diode
R659 N658 N659 10
D659 N659 0 diode
R660 N659 N660 10
D660 N660 0 diode
R661 N660 N661 10
D661 N661 0 diode
R662 N661 N662 10
D662 N662 0 diode
R663 N662 N663 10
D663 N663 0 diode
R664 N663 N664 10
D664 N664 0 diode
R665 N664 N665 10
D665 N665 0 diode
R666 N665 N666 10
D666 N666 0 diode
R667 N666 N667 10
D667 N667 0 diode
R668 N667 N668 10
D668 N668 0 diode
R669 N668 N669 10
D669 N669 0 diode
R670 N669 N670 10
D670 N670 0 diode
R671 N670 N671 10
D671 N671 0 diode
R672 N671 N672 10
D672 N672 0 diode
R673 N672 N673 10
D673 N673 0 diode
R674 N673 N674 10
D674 N674 0 diode
R675 N674 N675 10
D675 N675 0 diode
R676 N675 N676 10
D676 N676 0 diode
R677 N676 N677 10
D677 N677 0 diode
R678 N677 N678 10
D678 N678 0 diode
R679 N678 N679 10
D679 N679 0 diode
R680 N679 N680 10
D680 N680 0 diode
R681 N680 N681 10
D681 N681 0 diode
R682 N681 N682 10
D682 N682 0 diode
R683 N682 N683 10
D683 N683 0 diode
R684 N683 N684 10
D684 N684 0 diode
R685 N684 N685 10
D685 N685 0 diode
R686 N685 N686 10
D686 N686 0 diode
R687 N686 N687 10
D687 N687 0 diode
R688 N687 N688 10
D688 N688 0 diode
R689 N688 N689 10
D689 N689 0 diode
R690 N689 N690 10
D690 N690 0 diode
R691 N690 N691 10
D691 N691 0 diode
R692 N691 N692 10
D692 N692 0 diode
R693 N692 N693 10
D693 N693 0 diode
R694 N693 N694 10
D694 N694 0 diode
R695 N694 N695 10
D695 N695 0 diode
R696 N695 N696 10
D696 N696 0 diode
R697 N696 N697 10
D697 N697 0 diode
R698 N697 N698 10
D698 N698 0 diode
R699 N698 N699 10
D699 N699 0 diode
R700 N699 N700 10
D700 N700 0 diode
R701 N700 N701 10
D701 N701 0 diode
R702 N701 N702 10
D702 N702 0 diode
R703 N702 N703 10
D703 N703 0 diode
R704 N703 N704 10
D704 N704 0 diode
R705 N704 N705 10
D705 N705 0 diode
R706 N705 N706 10
D706 N706 0 diode
R707 N706 N707 10
D707 N707 0 diode
R708 N707 N708 10
D708 N708 0 diode
R709 N708 N709 10
D709 N709 0 diode
R710 N709 N710 10
D710 N710 0 diode
R711 N710 N711 10
D711 N711 0 diode
R712 N711 N712 10
D712 N712 0 diode
R713 N712 N713 10
D713 N713 0 diode
R714 N713 N714 10
D714 N714 0 diode
R715 N714 N715 10
D715 N715 0 diode
R716 N715 N716 10
D716 N716 0 diode
R717 N716 N717 10
D717 N717 0 diode
R718 N717 N718 10
D718 N718 0 diode
R719 N718 N719 10
D719 N719 0 diode
R720 N719 N720 10
D720 N720 0 diode
R721 N720 N721 10
D721 N721 0 diode
R722 N721 N722 10
D722 N722 0 diode
R723 N722 N723 10
D723 N723 0 diode
R724 N723 N724 10
D724 N724 0 diode
R725 N724 N725 10
D725 N725 0 diode
R726 N725 N726 10
D726 N726 0 diode
R727 N726 N727 10
D727 N727 0 diode
R728 N727 N728 10
D728 N728 0 diode
R729 N728 N729 10
D729 N729 0 diode
R730 N729 N730 10
D730 N730 0 diode
R731 N730 N731 10
D731 N731 0 diode
R732 N731 N732 10
D732 N732 0 diode
R733 N732 N733 10
D733 N733 0 diode
R734 N733 N734 10
D734 N734 0 diode
R735 N734 N735 10
D735 N735 0 diode
R736 N735 N736 10
D736 N736 0 diode
R737 N736 N737 10
D737 N737 0 diode
R738 N737 N738 10
D738 N738 0 diode
R739 N738 N739 10
D739 N739 0 diode
R740 N739 N740 10
D740 N740 0 diode
R741 N740 N741 10
D741 N741 0 diode
R742 N741 N742 10
D742 N742 0 diode
R743 N742 N743 10
D743 N743 0 diode
R744 N743 N744 10
D744 N744 0 diode
R745 N744 N745 10
D745 N745 0 diode
R746 N745 N746 10
D746 N746 0 diode
R747 N746 N747 10
D747 N747 0 diode
R748 N747 N748 10
D748 N748 0 diode
R749 N748 N749 10
D749 N749 0 diode
R750 N749 N750 10
D750 N750 0 diode
R751 N750 N751 10
D751 N751 0 diode
R752 N751 N752 10
D752 N752 0 diode
R753 N752 N753 10
D753 N753 0 diode
R754 N753 N754 10
D754 N754 0 diode
R755 N754 N755 10
D755 N755 0 diode
R756 N755 N756 10
D756 N756 0 diode
R757 N756 N757 10
D757 N757 0 diode
R758 N757 N758 10
D758 N758 0 diode
R759 N758 N759 10
D759 N759 0 diode
R760 N759 N760 10
D760 N760 0 diode
R761 N760 N761 10
D761 N761 0 diode
R762 N761 N762 10
D762 N762 0 diode
R763 N762 N763 10
D763 N763 0 diode
R764 N763 N764 10
D764 N764 0 diode
R765 N764 N765 10
D765 N765 0 diode
R766 N765 N766 10
D766 N766 0 diode
R767 N766 N767 10
D767 N767 0 diode
R768 N767 N768 10
D768 N768 0 diode
R769 N768 N769 10
D769 N769 0 diode
R770 N769 N770 10
D770 N770 0 diode
R771 N770 N771 10
D771 N771 0 diode
R772 N771 N772 10
D772 N772 0 diode
R773 N772 N773 10
D773 N773 0 diode
R774 N773 N774 10
D774 N774 0 diode
R775 N774 N775 10
D775 N775 0 diode
R776 N775 N776 10
D776 N776 0 diode
R777 N776 N777 10
D777 N777 0 diode
R778 N777 N778 10
D778 N778 0 diode
R779 N778 N779 10
D779 N779 0 diode
R780 N779 N780 10
D780 N780 0 diode
R781 N780 N781 10
D781 N781 0 diode
R782 N781 N782 10
D782 N782 0 diode
R783 N782 N783 10
D783 N783 0 diode
R784 N783 N784 10
D784 N784 0 diode
R785 N784 N785 10
D785 N785 0 diode
R786 N785 N786 10
D786 N786 0 diode
R787 N786 N787 10
D787 N787 0 diode
R788 N787 N788 10
D788 N788 0 diode
R789 N788 N789 10
D789 N789 0 diode
R790 N789 N790 10
D790 N790 0 diode
R791 N790 N791 10
D791 N791 0 diode
R792 N791 N792 10
D792 N792 0 diode
R793 N792 N793 10
D793 N793 0 diode
R794 N793 N794 10
D794 N794 0 diode
R795 N794 N795 10
D795 N795 0 diode
R796 N795 N796 10
D796 N796 0 diode
R797 N796 N797 10
D797 N797 0 diode
R798 N797 N798 10
D798 N798 0 diode
R799 N798 N799 10
D799 N799 0 diode
R800 N799 N800 10
D800 N800 0 diode
R801 N800 N801 10
D801 N801 0 diode
R802 N801 N802 10
D802 N802 0 diode
R803 N802 N803 10
D803 N803 0 diode
R804 N803 N804 10
D804 N804 0 diode
R805 N804 N805 10
D805 N805 0 diode
R806 N805 N806 10
D806 N806 0 diode
R807 N806 N807 10
D807 N807 0 diode
R808 N807 N808 10
D808 N808 0 diode
R809 N808 N809 10
D809 N809 0 diode
R810 N809 N810 10
D810 N810 0 diode
R811 N810 N811 10
D811 N811 0 diode
R812 N811 N812 10
D812 N812 0 diode
R813 N812 N813 10
D813 N813 0 diode
R814 N813 N814 10
D814 N814 0 diode
R815 N814 N815 10
D815 N815 0 diode
R816 N815 N816 10
D816 N816 0 diode
R817 N816 N817 10
D817 N817 0 diode
R818 N817 N818 10
D818 N818 0 diode
R819 N818 N819 10
D819 N819 0 diode
R820 N819 N820 10
D820 N820 0 diode
R821 N820 N821 10
D821 N821 0 diode
R822 N821 N822 10
D822 N822 0 diode
R823 N822 N823 10
D823 N823 0 diode
R824 N823 N824 10
D824 N824 0 diode
R825 N824 N825 10
D825 N825 0 diode
R826 N825 N826 10
D826 N826 0 diode
R827 N826 N827 10
D827 N827 0 diode
R828 N827 N828 10
D828 N828 0 diode
R829 N828 N829 10
D829 N829 0 diode
R830 N829 N830 10
D830 N830 0 diode
R831 N830 N831 10
D831 N831 0 diode
R832 N831 N832 10
D832 N832 0 diode
R833 N832 N833 10
D833 N833 0 diode
R834 N833 N834 10
D834 N834 0 diode
R835 N834 N835 10
D835 N835 0 diode
R836 N835 N836 10
D836 N836 0 diode
R837 N836 N837 10
D837 N837 0 diode
R838 N837 N838 10
D838 N838 0 diode
R839 N838 N839 10
D839 N839 0 diode
R840 N839 N840 10
D840 N840 0 diode
R841 N840 N841 10
D841 N841 0 diode
R842 N841 N842 10
D842 N842 0 diode
R843 N842 N843 10
D843 N843 0 diode
R844 N843 N844 10
D844 N844 0 diode
R845 N844 N845 10
D845 N845 0 diode
R846 N845 N846 10
D846 N846 0 diode
R847 N846 N847 10
D847 N847 0 diode
R848 N847 N848 10
D848 N848 0 diode
R849 N848 N849 10
D849 N849 0 diode
R850 N849 N850 10
D850 N850 0 diode
R851 N850 N851 10
D851 N851 0 diode
R852 N851 N852 10
D852 N852 0 diode
R853 N852 N853 10
D853 N853 0 diode
R854 N853 N854 10
D854 N854 0 diode
R855 N854 N855 10
D855 N855 0 diode
R856 N855 N856 10
D856 N856 0 diode
R857 N856 N857 10
D857 N857 0 diode
R858 N857 N858 10
D858 N858 0 diode
R859 N858 N859 10
D859 N859 0 diode
R860 N859 N860 10
D860 N860 0 diode
R861 N860 N861 10
D861 N861 0 diode
R862 N861 N862 10
D862 N862 0 diode
R863 N862 N863 10
D863 N863 0 diode
R864 N863 N864 10
D864 N864 0 diode
R865 N864 N865 10
D865 N865 0 diode
R866 N865 N866 10
D866 N866 0 diode
R867 N866 N867 10
D867 N867 0 diode
R868 N867 N868 10
D868 N868 0 diode
R869 N868 N869 10
D869 N869 0 diode
R870 N869 N870 10
D870 N870 0 diode
R871 N870 N871 10
D871 N871 0 diode
R872 N871 N872 10
D872 N872 0 diode
R873 N872 N873 10
D873 N873 0 diode
R874 N873 N874 10
D874 N874 0 diode
R875 N874 N875 10
D875 N875 0 diode
R876 N875 N876 10
D876 N876 0 diode
R877 N876 N877 10
D877 N877 0 diode
R878 N877 N878 10
D878 N878 0 diode
R879 N878 N879 10
D879 N879 0 diode
R880 N879 N880 10
D880 N880 0 diode
R881 N880 N881 10
D881 N881 0 diode
R882 N881 N882 10
D882 N882 0 diode
R883 N882 N883 10
D883 N883 0 diode
R884 N883 N884 10
D884 N884 0 diode
R885 N884 N885 10
D885 N885 0 diode
R886 N885 N886 10
D886 N886 0 diode
R887 N886 N887 10
D887 N887 0 diode
R888 N887 N888 10
D888 N888 0 diode
R889 N888 N889 10
D889 N889 0 diode
R890 N889 N890 10
D890 N890 0 diode
R891 N890 N891 10
D891 N891 0 diode
R892 N891 N892 10
D892 N892 0 diode
R893 N892 N893 10
D893 N893 0 diode
R894 N893 N894 10
D894 N894 0 diode
R895 N894 N895 10
D895 N895 0 diode
R896 N895 N896 10
D896 N896 0 diode
R897 N896 N897 10
D897 N897 0 diode
R898 N897 N898 10
D898 N898 0 diode
R899 N898 N899 10
D899 N899 0 diode
R900 N899 N900 10
D900 N900 0 diode
R901 N900 N901 10
D901 N901 0 diode
R902 N901 N902 10
D902 N902 0 diode
R903 N902 N903 10
D903 N903 0 diode
R904 N903 N904 10
D904 N904 0 diode
R905 N904 N905 10
D905 N905 0 diode
R906 N905 N906 10
D906 N906 0 diode
R907 N906 N907 10
D907 N907 0 diode
R908 N907 N908 10
D908 N908 0 diode
R909 N908 N909 10
D909 N909 0 diode
R910 N909 N910 10
D910 N910 0 diode
R911 N910 N911 10
D911 N911 0 diode
R912 N911 N912 10
D912 N912 0 diode
R913 N912 N913 10
D913 N913 0 diode
R914 N913 N914 10
D914 N914 0 diode
R915 N914 N915 10
D915 N915 0 diode
R916 N915 N916 10
D916 N916 0 diode
R917 N916 N917 10
D917 N917 0 diode
R918 N917 N918 10
D918 N918 0 diode
R919 N918 N919 10
D919 N919 0 diode
R920 N919 N920 10
D920 N920 0 diode
R921 N920 N921 10
D921 N921 0 diode
R922 N921 N922 10
D922 N922 0 diode
R923 N922 N923 10
D923 N923 0 diode
R924 N923 N924 10
D924 N924 0 diode
R925 N924 N925 10
D925 N925 0 diode
R926 N925 N926 10
D926 N926 0 diode
R927 N926 N927 10
D927 N927 0 diode
R928 N927 N928 10
D928 N928 0 diode
R929 N928 N929 10
D929 N929 0 diode
R930 N929 N930 10
D930 N930 0 diode
R931 N930 N931 10
D931 N931 0 diode
R932 N931 N932 10
D932 N932 0 diode
R933 N932 N933 10
D933 N933 0 diode
R934 N933 N934 10
D934 N934 0 diode
R935 N934 N935 10
D935 N935 0 diode
R936 N935 N936 10
D936 N936 0 diode
R937 N936 N937 10
D937 N937 0 diode
R938 N937 N938 10
D938 N938 0 diode
R939 N938 N939 10
D939 N939 0 diode
R940 N939 N940 10
D940 N940 0 diode
R941 N940 N941 10
D941 N941 0 diode
R942 N941 N942 10
D942 N942 0 diode
R943 N942 N943 10
D943 N943 0 diode
R944 N943 N944 10
D944 N944 0 diode
R945 N944 N945 10
D945 N945 0 diode
R946 N945 N946 10
D946 N946 0 diode
R947 N946 N947 10
D947 N947 0 diode
R948 N947 N948 10
D948 N948 0 diode
R949 N948 N949 10
D949 N949 0 diode
R950 N949 N950 10
D950 N950 0 diode
R951 N950 N951 10
D951 N951 0 diode
R952 N951 N952 10
D952 N952 0 diode
R953 N952 N953 10
D953 N953 0 diode
R954 N953 N954 10
D954 N954 0 diode
R955 N954 N955 10
D955 N955 0 diode
R956 N955 N956 10
D956 N956 0 diode
R957 N956 N957 10
D957 N957 0 diode
R958 N957 N958 10
D958 N958 0 diode
R959 N958 N959 10
D959 N959 0 diode
R960 N959 N960 10
D960 N960 0 diode
R961 N960 N961 10
D961 N961 0 diode
R962 N961 N962 10
D962 N962 0 diode
R963 N962 N963 10
D963 N963 0 diode
R964 N963 N964 10
D964 N964 0 diode
R965 N964 N965 10
D965 N965 0 diode
R966 N965 N966 10
D966 N966 0 diode
R967 N966 N967 10
D967 N967 0 diode
R968 N967 N968 10
D968 N968 0 diode
R969 N968 N969 10
D969 N969 0 diode
R970 N969 N970 10
D970 N970 0 diode
R971 N970 N971 10
D971 N971 0 diode
R972 N971 N972 10
D972 N972 0 diode
R973 N972 N973 10
D973 N973 0 diode
R974 N973 N974 10
D974 N974 0 diode
R975 N974 N975 10
D975 N975 0 diode
R976 N975 N976 10
D976 N976 0 diode
R977 N976 N977 10
D977 N977 0 diode
R978 N977 N978 10
D978 N978 0 diode
R979 N978 N979 10
D979 N979 0 diode
R980 N979 N980 10
D980 N980 0 diode
R981 N980 N981 10
D981 N981 0 diode
R982 N981 N982 10
D982 N982 0 diode
R983 N982 N983 10
D983 N983 0 diode
R984 N983 N984 10
D984 N984 0 diode
R985 N984 N985 10
D985 N985 0 diode
R986 N985 N986 10
D986 N986 0 diode
R987 N986 N987 10
D987 N987 0 diode
R988 N987 N988 10
D988 N988 0 diode
R989 N988 N989 10
D989 N989 0 diode
R990 N989 N990 10
D990 N990 0 diode
R991 N990 N991 10
D991 N991 0 diode
R992 N991 N992 10
D992 N992 0 diode
R993 N992 N993 10
D993 N993 0 diode
R994 N993 N994 10
D994 N994 0 diode
R995 N994 N995 10
D995 N995 0 diode
R996 N995 N996 10
D996 N996 0 diode
R997 N996 N997 10
D997 N997 0 diode
R998 N997 N998 10
D998 N998 0 diode
R999 N998 N999 10
D999 N999 0 diode
R1000 N999 N1000 10
D1000 N1000 0 diode
.op
.control                                    ; begin of control section
run                                         ; run the .tran command
print N50000
.endc 
.end