V1 0 1 10
R1 1 2 100
C1 2 3 0.001
L1 3 0 0.1
.tran 0.001 0.01