V1 0 RNODE 10
R1 RNODE 0 10
.tran 1e-3 1e-2