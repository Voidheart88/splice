* Test circuit with controlled sources

* Independent voltage source
Vin 1 0 10

* Resistors
R1 1 2 1000
R2 2 0 1000

* VCVS - Voltage-Controlled Voltage Source (E source)
* Output voltage = gain * (V(ctrl_pos) - V(ctrl_neg))
E1 3 0 2 0 2.0  ; V(3) = 2.0 * V(2)

* VCCS - Voltage-Controlled Current Source (G source)
* Output current = transconductance * (V(ctrl_pos) - V(ctrl_neg))
G1 3 4 2 0 0.01  ; I(3->4) = 0.01 * V(2)

* CCCS - Current-Controlled Current Source (F source)
* Output current = gain * I(ctrl_branch)
F1 5 6 V1 10.0  ; I(5->6) = 10.0 * I(V1)

* CCVS - Current-Controlled Voltage Source (H source)
* Output voltage = gain * I(ctrl_branch)
H1 7 0 V1 5.0  ; V(7) = 5.0 * I(V1)

* Analysis
.op
.end