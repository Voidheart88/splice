V1 0 1 5
R1 1 2 1000
C1 2 0 0.001
.tran 0.00001 10