V1 0 1 10
R1 1 2 100
L1 2 0 0.1
.tran 0.001 0.01