V1 0 1 STEP 0 10 0.5
L1 1 2 0.1
R1 2 0 10
.tran 0.1 10