V1 0 1 10
R1 1 2 1e3
C1 2 0 100e-9
.tran 1e-6 1e-3