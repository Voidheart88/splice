V1 0 1 SIN 0 10 1
.tran 1 10