V1 0 1 10
.tran 1 10