V1 0 1 10
L1 1 0 0.1
.tran 0.001 0.01