V1 1 0 DC 1
R1 1 2 1k
C1 2 0 1uF
.tran 1e-7 1e-3
.end
