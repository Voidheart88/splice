V1 0 1 10
R1 1 2 1000
C1 2 0 1000
.tran 1e-9 1e-6