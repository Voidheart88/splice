*Test*
.model diode D()
V1 N0 0 10
R1 N0 N1 10
D1 N1 0 diode
R2 N1 N2 10
D2 N2 0 diode
R3 N2 N3 10
D3 N3 0 diode
R4 N3 N4 10
D4 N4 0 diode
R5 N4 N5 10
D5 N5 0 diode
R6 N5 N6 10
D6 N6 0 diode
R7 N6 N7 10
D7 N7 0 diode
R8 N7 N8 10
D8 N8 0 diode
R9 N8 N9 10
D9 N9 0 diode
R10 N9 N10 10
D10 N10 0 diode
R11 N10 N11 10
D11 N11 0 diode
R12 N11 N12 10
D12 N12 0 diode
R13 N12 N13 10
D13 N13 0 diode
R14 N13 N14 10
D14 N14 0 diode
R15 N14 N15 10
D15 N15 0 diode
R16 N15 N16 10
D16 N16 0 diode
R17 N16 N17 10
D17 N17 0 diode
R18 N17 N18 10
D18 N18 0 diode
R19 N18 N19 10
D19 N19 0 diode
R20 N19 N20 10
D20 N20 0 diode
R21 N20 N21 10
D21 N21 0 diode
R22 N21 N22 10
D22 N22 0 diode
R23 N22 N23 10
D23 N23 0 diode
R24 N23 N24 10
D24 N24 0 diode
R25 N24 N25 10
D25 N25 0 diode
R26 N25 N26 10
D26 N26 0 diode
R27 N26 N27 10
D27 N27 0 diode
R28 N27 N28 10
D28 N28 0 diode
R29 N28 N29 10
D29 N29 0 diode
R30 N29 N30 10
D30 N30 0 diode
R31 N30 N31 10
D31 N31 0 diode
R32 N31 N32 10
D32 N32 0 diode
R33 N32 N33 10
D33 N33 0 diode
R34 N33 N34 10
D34 N34 0 diode
R35 N34 N35 10
D35 N35 0 diode
R36 N35 N36 10
D36 N36 0 diode
R37 N36 N37 10
D37 N37 0 diode
R38 N37 N38 10
D38 N38 0 diode
R39 N38 N39 10
D39 N39 0 diode
R40 N39 N40 10
D40 N40 0 diode
R41 N40 N41 10
D41 N41 0 diode
R42 N41 N42 10
D42 N42 0 diode
R43 N42 N43 10
D43 N43 0 diode
R44 N43 N44 10
D44 N44 0 diode
R45 N44 N45 10
D45 N45 0 diode
R46 N45 N46 10
D46 N46 0 diode
R47 N46 N47 10
D47 N47 0 diode
R48 N47 N48 10
D48 N48 0 diode
R49 N48 N49 10
D49 N49 0 diode
R50 N49 N50 10
D50 N50 0 diode
R51 N50 N51 10
D51 N51 0 diode
R52 N51 N52 10
D52 N52 0 diode
R53 N52 N53 10
D53 N53 0 diode
R54 N53 N54 10
D54 N54 0 diode
R55 N54 N55 10
D55 N55 0 diode
R56 N55 N56 10
D56 N56 0 diode
R57 N56 N57 10
D57 N57 0 diode
R58 N57 N58 10
D58 N58 0 diode
R59 N58 N59 10
D59 N59 0 diode
R60 N59 N60 10
D60 N60 0 diode
R61 N60 N61 10
D61 N61 0 diode
R62 N61 N62 10
D62 N62 0 diode
R63 N62 N63 10
D63 N63 0 diode
R64 N63 N64 10
D64 N64 0 diode
R65 N64 N65 10
D65 N65 0 diode
R66 N65 N66 10
D66 N66 0 diode
R67 N66 N67 10
D67 N67 0 diode
R68 N67 N68 10
D68 N68 0 diode
R69 N68 N69 10
D69 N69 0 diode
R70 N69 N70 10
D70 N70 0 diode
R71 N70 N71 10
D71 N71 0 diode
R72 N71 N72 10
D72 N72 0 diode
R73 N72 N73 10
D73 N73 0 diode
R74 N73 N74 10
D74 N74 0 diode
R75 N74 N75 10
D75 N75 0 diode
R76 N75 N76 10
D76 N76 0 diode
R77 N76 N77 10
D77 N77 0 diode
R78 N77 N78 10
D78 N78 0 diode
R79 N78 N79 10
D79 N79 0 diode
R80 N79 N80 10
D80 N80 0 diode
R81 N80 N81 10
D81 N81 0 diode
R82 N81 N82 10
D82 N82 0 diode
R83 N82 N83 10
D83 N83 0 diode
R84 N83 N84 10
D84 N84 0 diode
R85 N84 N85 10
D85 N85 0 diode
R86 N85 N86 10
D86 N86 0 diode
R87 N86 N87 10
D87 N87 0 diode
R88 N87 N88 10
D88 N88 0 diode
R89 N88 N89 10
D89 N89 0 diode
R90 N89 N90 10
D90 N90 0 diode
R91 N90 N91 10
D91 N91 0 diode
R92 N91 N92 10
D92 N92 0 diode
R93 N92 N93 10
D93 N93 0 diode
R94 N93 N94 10
D94 N94 0 diode
R95 N94 N95 10
D95 N95 0 diode
R96 N95 N96 10
D96 N96 0 diode
R97 N96 N97 10
D97 N97 0 diode
R98 N97 N98 10
D98 N98 0 diode
R99 N98 N99 10
D99 N99 0 diode
R100 N99 N100 10
D100 N100 0 diode
R101 N100 N101 10
D101 N101 0 diode
R102 N101 N102 10
D102 N102 0 diode
R103 N102 N103 10
D103 N103 0 diode
R104 N103 N104 10
D104 N104 0 diode
R105 N104 N105 10
D105 N105 0 diode
R106 N105 N106 10
D106 N106 0 diode
R107 N106 N107 10
D107 N107 0 diode
R108 N107 N108 10
D108 N108 0 diode
R109 N108 N109 10
D109 N109 0 diode
R110 N109 N110 10
D110 N110 0 diode
R111 N110 N111 10
D111 N111 0 diode
R112 N111 N112 10
D112 N112 0 diode
R113 N112 N113 10
D113 N113 0 diode
R114 N113 N114 10
D114 N114 0 diode
R115 N114 N115 10
D115 N115 0 diode
R116 N115 N116 10
D116 N116 0 diode
R117 N116 N117 10
D117 N117 0 diode
R118 N117 N118 10
D118 N118 0 diode
R119 N118 N119 10
D119 N119 0 diode
R120 N119 N120 10
D120 N120 0 diode
R121 N120 N121 10
D121 N121 0 diode
R122 N121 N122 10
D122 N122 0 diode
R123 N122 N123 10
D123 N123 0 diode
R124 N123 N124 10
D124 N124 0 diode
R125 N124 N125 10
D125 N125 0 diode
R126 N125 N126 10
D126 N126 0 diode
R127 N126 N127 10
D127 N127 0 diode
R128 N127 N128 10
D128 N128 0 diode
R129 N128 N129 10
D129 N129 0 diode
R130 N129 N130 10
D130 N130 0 diode
R131 N130 N131 10
D131 N131 0 diode
R132 N131 N132 10
D132 N132 0 diode
R133 N132 N133 10
D133 N133 0 diode
R134 N133 N134 10
D134 N134 0 diode
R135 N134 N135 10
D135 N135 0 diode
R136 N135 N136 10
D136 N136 0 diode
R137 N136 N137 10
D137 N137 0 diode
R138 N137 N138 10
D138 N138 0 diode
R139 N138 N139 10
D139 N139 0 diode
R140 N139 N140 10
D140 N140 0 diode
R141 N140 N141 10
D141 N141 0 diode
R142 N141 N142 10
D142 N142 0 diode
R143 N142 N143 10
D143 N143 0 diode
R144 N143 N144 10
D144 N144 0 diode
R145 N144 N145 10
D145 N145 0 diode
R146 N145 N146 10
D146 N146 0 diode
R147 N146 N147 10
D147 N147 0 diode
R148 N147 N148 10
D148 N148 0 diode
R149 N148 N149 10
D149 N149 0 diode
R150 N149 N150 10
D150 N150 0 diode
R151 N150 N151 10
D151 N151 0 diode
R152 N151 N152 10
D152 N152 0 diode
R153 N152 N153 10
D153 N153 0 diode
R154 N153 N154 10
D154 N154 0 diode
R155 N154 N155 10
D155 N155 0 diode
R156 N155 N156 10
D156 N156 0 diode
R157 N156 N157 10
D157 N157 0 diode
R158 N157 N158 10
D158 N158 0 diode
R159 N158 N159 10
D159 N159 0 diode
R160 N159 N160 10
D160 N160 0 diode
R161 N160 N161 10
D161 N161 0 diode
R162 N161 N162 10
D162 N162 0 diode
R163 N162 N163 10
D163 N163 0 diode
R164 N163 N164 10
D164 N164 0 diode
R165 N164 N165 10
D165 N165 0 diode
R166 N165 N166 10
D166 N166 0 diode
R167 N166 N167 10
D167 N167 0 diode
R168 N167 N168 10
D168 N168 0 diode
R169 N168 N169 10
D169 N169 0 diode
R170 N169 N170 10
D170 N170 0 diode
R171 N170 N171 10
D171 N171 0 diode
R172 N171 N172 10
D172 N172 0 diode
R173 N172 N173 10
D173 N173 0 diode
R174 N173 N174 10
D174 N174 0 diode
R175 N174 N175 10
D175 N175 0 diode
R176 N175 N176 10
D176 N176 0 diode
R177 N176 N177 10
D177 N177 0 diode
R178 N177 N178 10
D178 N178 0 diode
R179 N178 N179 10
D179 N179 0 diode
R180 N179 N180 10
D180 N180 0 diode
R181 N180 N181 10
D181 N181 0 diode
R182 N181 N182 10
D182 N182 0 diode
R183 N182 N183 10
D183 N183 0 diode
R184 N183 N184 10
D184 N184 0 diode
R185 N184 N185 10
D185 N185 0 diode
R186 N185 N186 10
D186 N186 0 diode
R187 N186 N187 10
D187 N187 0 diode
R188 N187 N188 10
D188 N188 0 diode
R189 N188 N189 10
D189 N189 0 diode
R190 N189 N190 10
D190 N190 0 diode
R191 N190 N191 10
D191 N191 0 diode
R192 N191 N192 10
D192 N192 0 diode
R193 N192 N193 10
D193 N193 0 diode
R194 N193 N194 10
D194 N194 0 diode
R195 N194 N195 10
D195 N195 0 diode
R196 N195 N196 10
D196 N196 0 diode
R197 N196 N197 10
D197 N197 0 diode
R198 N197 N198 10
D198 N198 0 diode
R199 N198 N199 10
D199 N199 0 diode
R200 N199 N200 10
D200 N200 0 diode
R201 N200 N201 10
D201 N201 0 diode
R202 N201 N202 10
D202 N202 0 diode
R203 N202 N203 10
D203 N203 0 diode
R204 N203 N204 10
D204 N204 0 diode
R205 N204 N205 10
D205 N205 0 diode
R206 N205 N206 10
D206 N206 0 diode
R207 N206 N207 10
D207 N207 0 diode
R208 N207 N208 10
D208 N208 0 diode
R209 N208 N209 10
D209 N209 0 diode
R210 N209 N210 10
D210 N210 0 diode
R211 N210 N211 10
D211 N211 0 diode
R212 N211 N212 10
D212 N212 0 diode
R213 N212 N213 10
D213 N213 0 diode
R214 N213 N214 10
D214 N214 0 diode
R215 N214 N215 10
D215 N215 0 diode
R216 N215 N216 10
D216 N216 0 diode
R217 N216 N217 10
D217 N217 0 diode
R218 N217 N218 10
D218 N218 0 diode
R219 N218 N219 10
D219 N219 0 diode
R220 N219 N220 10
D220 N220 0 diode
R221 N220 N221 10
D221 N221 0 diode
R222 N221 N222 10
D222 N222 0 diode
R223 N222 N223 10
D223 N223 0 diode
R224 N223 N224 10
D224 N224 0 diode
R225 N224 N225 10
D225 N225 0 diode
R226 N225 N226 10
D226 N226 0 diode
R227 N226 N227 10
D227 N227 0 diode
R228 N227 N228 10
D228 N228 0 diode
R229 N228 N229 10
D229 N229 0 diode
R230 N229 N230 10
D230 N230 0 diode
R231 N230 N231 10
D231 N231 0 diode
R232 N231 N232 10
D232 N232 0 diode
R233 N232 N233 10
D233 N233 0 diode
R234 N233 N234 10
D234 N234 0 diode
R235 N234 N235 10
D235 N235 0 diode
R236 N235 N236 10
D236 N236 0 diode
R237 N236 N237 10
D237 N237 0 diode
R238 N237 N238 10
D238 N238 0 diode
R239 N238 N239 10
D239 N239 0 diode
R240 N239 N240 10
D240 N240 0 diode
R241 N240 N241 10
D241 N241 0 diode
R242 N241 N242 10
D242 N242 0 diode
R243 N242 N243 10
D243 N243 0 diode
R244 N243 N244 10
D244 N244 0 diode
R245 N244 N245 10
D245 N245 0 diode
R246 N245 N246 10
D246 N246 0 diode
R247 N246 N247 10
D247 N247 0 diode
R248 N247 N248 10
D248 N248 0 diode
R249 N248 N249 10
D249 N249 0 diode
R250 N249 N250 10
D250 N250 0 diode
R251 N250 N251 10
D251 N251 0 diode
R252 N251 N252 10
D252 N252 0 diode
R253 N252 N253 10
D253 N253 0 diode
R254 N253 N254 10
D254 N254 0 diode
R255 N254 N255 10
D255 N255 0 diode
R256 N255 N256 10
D256 N256 0 diode
R257 N256 N257 10
D257 N257 0 diode
R258 N257 N258 10
D258 N258 0 diode
R259 N258 N259 10
D259 N259 0 diode
R260 N259 N260 10
D260 N260 0 diode
R261 N260 N261 10
D261 N261 0 diode
R262 N261 N262 10
D262 N262 0 diode
R263 N262 N263 10
D263 N263 0 diode
R264 N263 N264 10
D264 N264 0 diode
R265 N264 N265 10
D265 N265 0 diode
R266 N265 N266 10
D266 N266 0 diode
R267 N266 N267 10
D267 N267 0 diode
R268 N267 N268 10
D268 N268 0 diode
R269 N268 N269 10
D269 N269 0 diode
R270 N269 N270 10
D270 N270 0 diode
R271 N270 N271 10
D271 N271 0 diode
R272 N271 N272 10
D272 N272 0 diode
R273 N272 N273 10
D273 N273 0 diode
R274 N273 N274 10
D274 N274 0 diode
R275 N274 N275 10
D275 N275 0 diode
R276 N275 N276 10
D276 N276 0 diode
R277 N276 N277 10
D277 N277 0 diode
R278 N277 N278 10
D278 N278 0 diode
R279 N278 N279 10
D279 N279 0 diode
R280 N279 N280 10
D280 N280 0 diode
R281 N280 N281 10
D281 N281 0 diode
R282 N281 N282 10
D282 N282 0 diode
R283 N282 N283 10
D283 N283 0 diode
R284 N283 N284 10
D284 N284 0 diode
R285 N284 N285 10
D285 N285 0 diode
R286 N285 N286 10
D286 N286 0 diode
R287 N286 N287 10
D287 N287 0 diode
R288 N287 N288 10
D288 N288 0 diode
R289 N288 N289 10
D289 N289 0 diode
R290 N289 N290 10
D290 N290 0 diode
R291 N290 N291 10
D291 N291 0 diode
R292 N291 N292 10
D292 N292 0 diode
R293 N292 N293 10
D293 N293 0 diode
R294 N293 N294 10
D294 N294 0 diode
R295 N294 N295 10
D295 N295 0 diode
R296 N295 N296 10
D296 N296 0 diode
R297 N296 N297 10
D297 N297 0 diode
R298 N297 N298 10
D298 N298 0 diode
R299 N298 N299 10
D299 N299 0 diode
R300 N299 N300 10
D300 N300 0 diode
R301 N300 N301 10
D301 N301 0 diode
R302 N301 N302 10
D302 N302 0 diode
R303 N302 N303 10
D303 N303 0 diode
R304 N303 N304 10
D304 N304 0 diode
R305 N304 N305 10
D305 N305 0 diode
R306 N305 N306 10
D306 N306 0 diode
R307 N306 N307 10
D307 N307 0 diode
R308 N307 N308 10
D308 N308 0 diode
R309 N308 N309 10
D309 N309 0 diode
R310 N309 N310 10
D310 N310 0 diode
R311 N310 N311 10
D311 N311 0 diode
R312 N311 N312 10
D312 N312 0 diode
R313 N312 N313 10
D313 N313 0 diode
R314 N313 N314 10
D314 N314 0 diode
R315 N314 N315 10
D315 N315 0 diode
R316 N315 N316 10
D316 N316 0 diode
R317 N316 N317 10
D317 N317 0 diode
R318 N317 N318 10
D318 N318 0 diode
R319 N318 N319 10
D319 N319 0 diode
R320 N319 N320 10
D320 N320 0 diode
R321 N320 N321 10
D321 N321 0 diode
R322 N321 N322 10
D322 N322 0 diode
R323 N322 N323 10
D323 N323 0 diode
R324 N323 N324 10
D324 N324 0 diode
R325 N324 N325 10
D325 N325 0 diode
R326 N325 N326 10
D326 N326 0 diode
R327 N326 N327 10
D327 N327 0 diode
R328 N327 N328 10
D328 N328 0 diode
R329 N328 N329 10
D329 N329 0 diode
R330 N329 N330 10
D330 N330 0 diode
R331 N330 N331 10
D331 N331 0 diode
R332 N331 N332 10
D332 N332 0 diode
R333 N332 N333 10
D333 N333 0 diode
R334 N333 N334 10
D334 N334 0 diode
R335 N334 N335 10
D335 N335 0 diode
R336 N335 N336 10
D336 N336 0 diode
R337 N336 N337 10
D337 N337 0 diode
R338 N337 N338 10
D338 N338 0 diode
R339 N338 N339 10
D339 N339 0 diode
R340 N339 N340 10
D340 N340 0 diode
R341 N340 N341 10
D341 N341 0 diode
R342 N341 N342 10
D342 N342 0 diode
R343 N342 N343 10
D343 N343 0 diode
R344 N343 N344 10
D344 N344 0 diode
R345 N344 N345 10
D345 N345 0 diode
R346 N345 N346 10
D346 N346 0 diode
R347 N346 N347 10
D347 N347 0 diode
R348 N347 N348 10
D348 N348 0 diode
R349 N348 N349 10
D349 N349 0 diode
R350 N349 N350 10
D350 N350 0 diode
R351 N350 N351 10
D351 N351 0 diode
R352 N351 N352 10
D352 N352 0 diode
R353 N352 N353 10
D353 N353 0 diode
R354 N353 N354 10
D354 N354 0 diode
R355 N354 N355 10
D355 N355 0 diode
R356 N355 N356 10
D356 N356 0 diode
R357 N356 N357 10
D357 N357 0 diode
R358 N357 N358 10
D358 N358 0 diode
R359 N358 N359 10
D359 N359 0 diode
R360 N359 N360 10
D360 N360 0 diode
R361 N360 N361 10
D361 N361 0 diode
R362 N361 N362 10
D362 N362 0 diode
R363 N362 N363 10
D363 N363 0 diode
R364 N363 N364 10
D364 N364 0 diode
R365 N364 N365 10
D365 N365 0 diode
R366 N365 N366 10
D366 N366 0 diode
R367 N366 N367 10
D367 N367 0 diode
R368 N367 N368 10
D368 N368 0 diode
R369 N368 N369 10
D369 N369 0 diode
R370 N369 N370 10
D370 N370 0 diode
R371 N370 N371 10
D371 N371 0 diode
R372 N371 N372 10
D372 N372 0 diode
R373 N372 N373 10
D373 N373 0 diode
R374 N373 N374 10
D374 N374 0 diode
R375 N374 N375 10
D375 N375 0 diode
R376 N375 N376 10
D376 N376 0 diode
R377 N376 N377 10
D377 N377 0 diode
R378 N377 N378 10
D378 N378 0 diode
R379 N378 N379 10
D379 N379 0 diode
R380 N379 N380 10
D380 N380 0 diode
R381 N380 N381 10
D381 N381 0 diode
R382 N381 N382 10
D382 N382 0 diode
R383 N382 N383 10
D383 N383 0 diode
R384 N383 N384 10
D384 N384 0 diode
R385 N384 N385 10
D385 N385 0 diode
R386 N385 N386 10
D386 N386 0 diode
R387 N386 N387 10
D387 N387 0 diode
R388 N387 N388 10
D388 N388 0 diode
R389 N388 N389 10
D389 N389 0 diode
R390 N389 N390 10
D390 N390 0 diode
R391 N390 N391 10
D391 N391 0 diode
R392 N391 N392 10
D392 N392 0 diode
R393 N392 N393 10
D393 N393 0 diode
R394 N393 N394 10
D394 N394 0 diode
R395 N394 N395 10
D395 N395 0 diode
R396 N395 N396 10
D396 N396 0 diode
R397 N396 N397 10
D397 N397 0 diode
R398 N397 N398 10
D398 N398 0 diode
R399 N398 N399 10
D399 N399 0 diode
R400 N399 N400 10
D400 N400 0 diode
R401 N400 N401 10
D401 N401 0 diode
R402 N401 N402 10
D402 N402 0 diode
R403 N402 N403 10
D403 N403 0 diode
R404 N403 N404 10
D404 N404 0 diode
R405 N404 N405 10
D405 N405 0 diode
R406 N405 N406 10
D406 N406 0 diode
R407 N406 N407 10
D407 N407 0 diode
R408 N407 N408 10
D408 N408 0 diode
R409 N408 N409 10
D409 N409 0 diode
R410 N409 N410 10
D410 N410 0 diode
R411 N410 N411 10
D411 N411 0 diode
R412 N411 N412 10
D412 N412 0 diode
R413 N412 N413 10
D413 N413 0 diode
R414 N413 N414 10
D414 N414 0 diode
R415 N414 N415 10
D415 N415 0 diode
R416 N415 N416 10
D416 N416 0 diode
R417 N416 N417 10
D417 N417 0 diode
R418 N417 N418 10
D418 N418 0 diode
R419 N418 N419 10
D419 N419 0 diode
R420 N419 N420 10
D420 N420 0 diode
R421 N420 N421 10
D421 N421 0 diode
R422 N421 N422 10
D422 N422 0 diode
R423 N422 N423 10
D423 N423 0 diode
R424 N423 N424 10
D424 N424 0 diode
R425 N424 N425 10
D425 N425 0 diode
R426 N425 N426 10
D426 N426 0 diode
R427 N426 N427 10
D427 N427 0 diode
R428 N427 N428 10
D428 N428 0 diode
R429 N428 N429 10
D429 N429 0 diode
R430 N429 N430 10
D430 N430 0 diode
R431 N430 N431 10
D431 N431 0 diode
R432 N431 N432 10
D432 N432 0 diode
R433 N432 N433 10
D433 N433 0 diode
R434 N433 N434 10
D434 N434 0 diode
R435 N434 N435 10
D435 N435 0 diode
R436 N435 N436 10
D436 N436 0 diode
R437 N436 N437 10
D437 N437 0 diode
R438 N437 N438 10
D438 N438 0 diode
R439 N438 N439 10
D439 N439 0 diode
R440 N439 N440 10
D440 N440 0 diode
R441 N440 N441 10
D441 N441 0 diode
R442 N441 N442 10
D442 N442 0 diode
R443 N442 N443 10
D443 N443 0 diode
R444 N443 N444 10
D444 N444 0 diode
R445 N444 N445 10
D445 N445 0 diode
R446 N445 N446 10
D446 N446 0 diode
R447 N446 N447 10
D447 N447 0 diode
R448 N447 N448 10
D448 N448 0 diode
R449 N448 N449 10
D449 N449 0 diode
R450 N449 N450 10
D450 N450 0 diode
R451 N450 N451 10
D451 N451 0 diode
R452 N451 N452 10
D452 N452 0 diode
R453 N452 N453 10
D453 N453 0 diode
R454 N453 N454 10
D454 N454 0 diode
R455 N454 N455 10
D455 N455 0 diode
R456 N455 N456 10
D456 N456 0 diode
R457 N456 N457 10
D457 N457 0 diode
R458 N457 N458 10
D458 N458 0 diode
R459 N458 N459 10
D459 N459 0 diode
R460 N459 N460 10
D460 N460 0 diode
R461 N460 N461 10
D461 N461 0 diode
R462 N461 N462 10
D462 N462 0 diode
R463 N462 N463 10
D463 N463 0 diode
R464 N463 N464 10
D464 N464 0 diode
R465 N464 N465 10
D465 N465 0 diode
R466 N465 N466 10
D466 N466 0 diode
R467 N466 N467 10
D467 N467 0 diode
R468 N467 N468 10
D468 N468 0 diode
R469 N468 N469 10
D469 N469 0 diode
R470 N469 N470 10
D470 N470 0 diode
R471 N470 N471 10
D471 N471 0 diode
R472 N471 N472 10
D472 N472 0 diode
R473 N472 N473 10
D473 N473 0 diode
R474 N473 N474 10
D474 N474 0 diode
R475 N474 N475 10
D475 N475 0 diode
R476 N475 N476 10
D476 N476 0 diode
R477 N476 N477 10
D477 N477 0 diode
R478 N477 N478 10
D478 N478 0 diode
R479 N478 N479 10
D479 N479 0 diode
R480 N479 N480 10
D480 N480 0 diode
R481 N480 N481 10
D481 N481 0 diode
R482 N481 N482 10
D482 N482 0 diode
R483 N482 N483 10
D483 N483 0 diode
R484 N483 N484 10
D484 N484 0 diode
R485 N484 N485 10
D485 N485 0 diode
R486 N485 N486 10
D486 N486 0 diode
R487 N486 N487 10
D487 N487 0 diode
R488 N487 N488 10
D488 N488 0 diode
R489 N488 N489 10
D489 N489 0 diode
R490 N489 N490 10
D490 N490 0 diode
R491 N490 N491 10
D491 N491 0 diode
R492 N491 N492 10
D492 N492 0 diode
R493 N492 N493 10
D493 N493 0 diode
R494 N493 N494 10
D494 N494 0 diode
R495 N494 N495 10
D495 N495 0 diode
R496 N495 N496 10
D496 N496 0 diode
R497 N496 N497 10
D497 N497 0 diode
R498 N497 N498 10
D498 N498 0 diode
R499 N498 N499 10
D499 N499 0 diode
R500 N499 N500 10
D500 N500 0 diode
R501 N500 N501 10
D501 N501 0 diode
R502 N501 N502 10
D502 N502 0 diode
R503 N502 N503 10
D503 N503 0 diode
R504 N503 N504 10
D504 N504 0 diode
R505 N504 N505 10
D505 N505 0 diode
R506 N505 N506 10
D506 N506 0 diode
R507 N506 N507 10
D507 N507 0 diode
R508 N507 N508 10
D508 N508 0 diode
R509 N508 N509 10
D509 N509 0 diode
R510 N509 N510 10
D510 N510 0 diode
R511 N510 N511 10
D511 N511 0 diode
R512 N511 N512 10
D512 N512 0 diode
R513 N512 N513 10
D513 N513 0 diode
R514 N513 N514 10
D514 N514 0 diode
R515 N514 N515 10
D515 N515 0 diode
R516 N515 N516 10
D516 N516 0 diode
R517 N516 N517 10
D517 N517 0 diode
R518 N517 N518 10
D518 N518 0 diode
R519 N518 N519 10
D519 N519 0 diode
R520 N519 N520 10
D520 N520 0 diode
R521 N520 N521 10
D521 N521 0 diode
R522 N521 N522 10
D522 N522 0 diode
R523 N522 N523 10
D523 N523 0 diode
R524 N523 N524 10
D524 N524 0 diode
R525 N524 N525 10
D525 N525 0 diode
R526 N525 N526 10
D526 N526 0 diode
R527 N526 N527 10
D527 N527 0 diode
R528 N527 N528 10
D528 N528 0 diode
R529 N528 N529 10
D529 N529 0 diode
R530 N529 N530 10
D530 N530 0 diode
R531 N530 N531 10
D531 N531 0 diode
R532 N531 N532 10
D532 N532 0 diode
R533 N532 N533 10
D533 N533 0 diode
R534 N533 N534 10
D534 N534 0 diode
R535 N534 N535 10
D535 N535 0 diode
R536 N535 N536 10
D536 N536 0 diode
R537 N536 N537 10
D537 N537 0 diode
R538 N537 N538 10
D538 N538 0 diode
R539 N538 N539 10
D539 N539 0 diode
R540 N539 N540 10
D540 N540 0 diode
R541 N540 N541 10
D541 N541 0 diode
R542 N541 N542 10
D542 N542 0 diode
R543 N542 N543 10
D543 N543 0 diode
R544 N543 N544 10
D544 N544 0 diode
R545 N544 N545 10
D545 N545 0 diode
R546 N545 N546 10
D546 N546 0 diode
R547 N546 N547 10
D547 N547 0 diode
R548 N547 N548 10
D548 N548 0 diode
R549 N548 N549 10
D549 N549 0 diode
R550 N549 N550 10
D550 N550 0 diode
R551 N550 N551 10
D551 N551 0 diode
R552 N551 N552 10
D552 N552 0 diode
R553 N552 N553 10
D553 N553 0 diode
R554 N553 N554 10
D554 N554 0 diode
R555 N554 N555 10
D555 N555 0 diode
R556 N555 N556 10
D556 N556 0 diode
R557 N556 N557 10
D557 N557 0 diode
R558 N557 N558 10
D558 N558 0 diode
R559 N558 N559 10
D559 N559 0 diode
R560 N559 N560 10
D560 N560 0 diode
R561 N560 N561 10
D561 N561 0 diode
R562 N561 N562 10
D562 N562 0 diode
R563 N562 N563 10
D563 N563 0 diode
R564 N563 N564 10
D564 N564 0 diode
R565 N564 N565 10
D565 N565 0 diode
R566 N565 N566 10
D566 N566 0 diode
R567 N566 N567 10
D567 N567 0 diode
R568 N567 N568 10
D568 N568 0 diode
R569 N568 N569 10
D569 N569 0 diode
R570 N569 N570 10
D570 N570 0 diode
R571 N570 N571 10
D571 N571 0 diode
R572 N571 N572 10
D572 N572 0 diode
R573 N572 N573 10
D573 N573 0 diode
R574 N573 N574 10
D574 N574 0 diode
R575 N574 N575 10
D575 N575 0 diode
R576 N575 N576 10
D576 N576 0 diode
R577 N576 N577 10
D577 N577 0 diode
R578 N577 N578 10
D578 N578 0 diode
R579 N578 N579 10
D579 N579 0 diode
R580 N579 N580 10
D580 N580 0 diode
R581 N580 N581 10
D581 N581 0 diode
R582 N581 N582 10
D582 N582 0 diode
R583 N582 N583 10
D583 N583 0 diode
R584 N583 N584 10
D584 N584 0 diode
R585 N584 N585 10
D585 N585 0 diode
R586 N585 N586 10
D586 N586 0 diode
R587 N586 N587 10
D587 N587 0 diode
R588 N587 N588 10
D588 N588 0 diode
R589 N588 N589 10
D589 N589 0 diode
R590 N589 N590 10
D590 N590 0 diode
R591 N590 N591 10
D591 N591 0 diode
R592 N591 N592 10
D592 N592 0 diode
R593 N592 N593 10
D593 N593 0 diode
R594 N593 N594 10
D594 N594 0 diode
R595 N594 N595 10
D595 N595 0 diode
R596 N595 N596 10
D596 N596 0 diode
R597 N596 N597 10
D597 N597 0 diode
R598 N597 N598 10
D598 N598 0 diode
R599 N598 N599 10
D599 N599 0 diode
R600 N599 N600 10
D600 N600 0 diode
R601 N600 N601 10
D601 N601 0 diode
R602 N601 N602 10
D602 N602 0 diode
R603 N602 N603 10
D603 N603 0 diode
R604 N603 N604 10
D604 N604 0 diode
R605 N604 N605 10
D605 N605 0 diode
R606 N605 N606 10
D606 N606 0 diode
R607 N606 N607 10
D607 N607 0 diode
R608 N607 N608 10
D608 N608 0 diode
R609 N608 N609 10
D609 N609 0 diode
R610 N609 N610 10
D610 N610 0 diode
R611 N610 N611 10
D611 N611 0 diode
R612 N611 N612 10
D612 N612 0 diode
R613 N612 N613 10
D613 N613 0 diode
R614 N613 N614 10
D614 N614 0 diode
R615 N614 N615 10
D615 N615 0 diode
R616 N615 N616 10
D616 N616 0 diode
R617 N616 N617 10
D617 N617 0 diode
R618 N617 N618 10
D618 N618 0 diode
R619 N618 N619 10
D619 N619 0 diode
R620 N619 N620 10
D620 N620 0 diode
R621 N620 N621 10
D621 N621 0 diode
R622 N621 N622 10
D622 N622 0 diode
R623 N622 N623 10
D623 N623 0 diode
R624 N623 N624 10
D624 N624 0 diode
R625 N624 N625 10
D625 N625 0 diode
R626 N625 N626 10
D626 N626 0 diode
R627 N626 N627 10
D627 N627 0 diode
R628 N627 N628 10
D628 N628 0 diode
R629 N628 N629 10
D629 N629 0 diode
R630 N629 N630 10
D630 N630 0 diode
R631 N630 N631 10
D631 N631 0 diode
R632 N631 N632 10
D632 N632 0 diode
R633 N632 N633 10
D633 N633 0 diode
R634 N633 N634 10
D634 N634 0 diode
R635 N634 N635 10
D635 N635 0 diode
R636 N635 N636 10
D636 N636 0 diode
R637 N636 N637 10
D637 N637 0 diode
R638 N637 N638 10
D638 N638 0 diode
R639 N638 N639 10
D639 N639 0 diode
R640 N639 N640 10
D640 N640 0 diode
R641 N640 N641 10
D641 N641 0 diode
R642 N641 N642 10
D642 N642 0 diode
R643 N642 N643 10
D643 N643 0 diode
R644 N643 N644 10
D644 N644 0 diode
R645 N644 N645 10
D645 N645 0 diode
R646 N645 N646 10
D646 N646 0 diode
R647 N646 N647 10
D647 N647 0 diode
R648 N647 N648 10
D648 N648 0 diode
R649 N648 N649 10
D649 N649 0 diode
R650 N649 N650 10
D650 N650 0 diode
R651 N650 N651 10
D651 N651 0 diode
R652 N651 N652 10
D652 N652 0 diode
R653 N652 N653 10
D653 N653 0 diode
R654 N653 N654 10
D654 N654 0 diode
R655 N654 N655 10
D655 N655 0 diode
R656 N655 N656 10
D656 N656 0 diode
R657 N656 N657 10
D657 N657 0 diode
R658 N657 N658 10
D658 N658 0 diode
R659 N658 N659 10
D659 N659 0 diode
R660 N659 N660 10
D660 N660 0 diode
R661 N660 N661 10
D661 N661 0 diode
R662 N661 N662 10
D662 N662 0 diode
R663 N662 N663 10
D663 N663 0 diode
R664 N663 N664 10
D664 N664 0 diode
R665 N664 N665 10
D665 N665 0 diode
R666 N665 N666 10
D666 N666 0 diode
R667 N666 N667 10
D667 N667 0 diode
R668 N667 N668 10
D668 N668 0 diode
R669 N668 N669 10
D669 N669 0 diode
R670 N669 N670 10
D670 N670 0 diode
R671 N670 N671 10
D671 N671 0 diode
R672 N671 N672 10
D672 N672 0 diode
R673 N672 N673 10
D673 N673 0 diode
R674 N673 N674 10
D674 N674 0 diode
R675 N674 N675 10
D675 N675 0 diode
R676 N675 N676 10
D676 N676 0 diode
R677 N676 N677 10
D677 N677 0 diode
R678 N677 N678 10
D678 N678 0 diode
R679 N678 N679 10
D679 N679 0 diode
R680 N679 N680 10
D680 N680 0 diode
R681 N680 N681 10
D681 N681 0 diode
R682 N681 N682 10
D682 N682 0 diode
R683 N682 N683 10
D683 N683 0 diode
R684 N683 N684 10
D684 N684 0 diode
R685 N684 N685 10
D685 N685 0 diode
R686 N685 N686 10
D686 N686 0 diode
R687 N686 N687 10
D687 N687 0 diode
R688 N687 N688 10
D688 N688 0 diode
R689 N688 N689 10
D689 N689 0 diode
R690 N689 N690 10
D690 N690 0 diode
R691 N690 N691 10
D691 N691 0 diode
R692 N691 N692 10
D692 N692 0 diode
R693 N692 N693 10
D693 N693 0 diode
R694 N693 N694 10
D694 N694 0 diode
R695 N694 N695 10
D695 N695 0 diode
R696 N695 N696 10
D696 N696 0 diode
R697 N696 N697 10
D697 N697 0 diode
R698 N697 N698 10
D698 N698 0 diode
R699 N698 N699 10
D699 N699 0 diode
R700 N699 N700 10
D700 N700 0 diode
R701 N700 N701 10
D701 N701 0 diode
R702 N701 N702 10
D702 N702 0 diode
R703 N702 N703 10
D703 N703 0 diode
R704 N703 N704 10
D704 N704 0 diode
R705 N704 N705 10
D705 N705 0 diode
R706 N705 N706 10
D706 N706 0 diode
R707 N706 N707 10
D707 N707 0 diode
R708 N707 N708 10
D708 N708 0 diode
R709 N708 N709 10
D709 N709 0 diode
R710 N709 N710 10
D710 N710 0 diode
R711 N710 N711 10
D711 N711 0 diode
R712 N711 N712 10
D712 N712 0 diode
R713 N712 N713 10
D713 N713 0 diode
R714 N713 N714 10
D714 N714 0 diode
R715 N714 N715 10
D715 N715 0 diode
R716 N715 N716 10
D716 N716 0 diode
R717 N716 N717 10
D717 N717 0 diode
R718 N717 N718 10
D718 N718 0 diode
R719 N718 N719 10
D719 N719 0 diode
R720 N719 N720 10
D720 N720 0 diode
R721 N720 N721 10
D721 N721 0 diode
R722 N721 N722 10
D722 N722 0 diode
R723 N722 N723 10
D723 N723 0 diode
R724 N723 N724 10
D724 N724 0 diode
R725 N724 N725 10
D725 N725 0 diode
R726 N725 N726 10
D726 N726 0 diode
R727 N726 N727 10
D727 N727 0 diode
R728 N727 N728 10
D728 N728 0 diode
R729 N728 N729 10
D729 N729 0 diode
R730 N729 N730 10
D730 N730 0 diode
R731 N730 N731 10
D731 N731 0 diode
R732 N731 N732 10
D732 N732 0 diode
R733 N732 N733 10
D733 N733 0 diode
R734 N733 N734 10
D734 N734 0 diode
R735 N734 N735 10
D735 N735 0 diode
R736 N735 N736 10
D736 N736 0 diode
R737 N736 N737 10
D737 N737 0 diode
R738 N737 N738 10
D738 N738 0 diode
R739 N738 N739 10
D739 N739 0 diode
R740 N739 N740 10
D740 N740 0 diode
R741 N740 N741 10
D741 N741 0 diode
R742 N741 N742 10
D742 N742 0 diode
R743 N742 N743 10
D743 N743 0 diode
R744 N743 N744 10
D744 N744 0 diode
R745 N744 N745 10
D745 N745 0 diode
R746 N745 N746 10
D746 N746 0 diode
R747 N746 N747 10
D747 N747 0 diode
R748 N747 N748 10
D748 N748 0 diode
R749 N748 N749 10
D749 N749 0 diode
R750 N749 N750 10
D750 N750 0 diode
R751 N750 N751 10
D751 N751 0 diode
R752 N751 N752 10
D752 N752 0 diode
R753 N752 N753 10
D753 N753 0 diode
R754 N753 N754 10
D754 N754 0 diode
R755 N754 N755 10
D755 N755 0 diode
R756 N755 N756 10
D756 N756 0 diode
R757 N756 N757 10
D757 N757 0 diode
R758 N757 N758 10
D758 N758 0 diode
R759 N758 N759 10
D759 N759 0 diode
R760 N759 N760 10
D760 N760 0 diode
R761 N760 N761 10
D761 N761 0 diode
R762 N761 N762 10
D762 N762 0 diode
R763 N762 N763 10
D763 N763 0 diode
R764 N763 N764 10
D764 N764 0 diode
R765 N764 N765 10
D765 N765 0 diode
R766 N765 N766 10
D766 N766 0 diode
R767 N766 N767 10
D767 N767 0 diode
R768 N767 N768 10
D768 N768 0 diode
R769 N768 N769 10
D769 N769 0 diode
R770 N769 N770 10
D770 N770 0 diode
R771 N770 N771 10
D771 N771 0 diode
R772 N771 N772 10
D772 N772 0 diode
R773 N772 N773 10
D773 N773 0 diode
R774 N773 N774 10
D774 N774 0 diode
R775 N774 N775 10
D775 N775 0 diode
R776 N775 N776 10
D776 N776 0 diode
R777 N776 N777 10
D777 N777 0 diode
R778 N777 N778 10
D778 N778 0 diode
R779 N778 N779 10
D779 N779 0 diode
R780 N779 N780 10
D780 N780 0 diode
R781 N780 N781 10
D781 N781 0 diode
R782 N781 N782 10
D782 N782 0 diode
R783 N782 N783 10
D783 N783 0 diode
R784 N783 N784 10
D784 N784 0 diode
R785 N784 N785 10
D785 N785 0 diode
R786 N785 N786 10
D786 N786 0 diode
R787 N786 N787 10
D787 N787 0 diode
R788 N787 N788 10
D788 N788 0 diode
R789 N788 N789 10
D789 N789 0 diode
R790 N789 N790 10
D790 N790 0 diode
R791 N790 N791 10
D791 N791 0 diode
R792 N791 N792 10
D792 N792 0 diode
R793 N792 N793 10
D793 N793 0 diode
R794 N793 N794 10
D794 N794 0 diode
R795 N794 N795 10
D795 N795 0 diode
R796 N795 N796 10
D796 N796 0 diode
R797 N796 N797 10
D797 N797 0 diode
R798 N797 N798 10
D798 N798 0 diode
R799 N798 N799 10
D799 N799 0 diode
R800 N799 N800 10
D800 N800 0 diode
R801 N800 N801 10
D801 N801 0 diode
R802 N801 N802 10
D802 N802 0 diode
R803 N802 N803 10
D803 N803 0 diode
R804 N803 N804 10
D804 N804 0 diode
R805 N804 N805 10
D805 N805 0 diode
R806 N805 N806 10
D806 N806 0 diode
R807 N806 N807 10
D807 N807 0 diode
R808 N807 N808 10
D808 N808 0 diode
R809 N808 N809 10
D809 N809 0 diode
R810 N809 N810 10
D810 N810 0 diode
R811 N810 N811 10
D811 N811 0 diode
R812 N811 N812 10
D812 N812 0 diode
R813 N812 N813 10
D813 N813 0 diode
R814 N813 N814 10
D814 N814 0 diode
R815 N814 N815 10
D815 N815 0 diode
R816 N815 N816 10
D816 N816 0 diode
R817 N816 N817 10
D817 N817 0 diode
R818 N817 N818 10
D818 N818 0 diode
R819 N818 N819 10
D819 N819 0 diode
R820 N819 N820 10
D820 N820 0 diode
R821 N820 N821 10
D821 N821 0 diode
R822 N821 N822 10
D822 N822 0 diode
R823 N822 N823 10
D823 N823 0 diode
R824 N823 N824 10
D824 N824 0 diode
R825 N824 N825 10
D825 N825 0 diode
R826 N825 N826 10
D826 N826 0 diode
R827 N826 N827 10
D827 N827 0 diode
R828 N827 N828 10
D828 N828 0 diode
R829 N828 N829 10
D829 N829 0 diode
R830 N829 N830 10
D830 N830 0 diode
R831 N830 N831 10
D831 N831 0 diode
R832 N831 N832 10
D832 N832 0 diode
R833 N832 N833 10
D833 N833 0 diode
R834 N833 N834 10
D834 N834 0 diode
R835 N834 N835 10
D835 N835 0 diode
R836 N835 N836 10
D836 N836 0 diode
R837 N836 N837 10
D837 N837 0 diode
R838 N837 N838 10
D838 N838 0 diode
R839 N838 N839 10
D839 N839 0 diode
R840 N839 N840 10
D840 N840 0 diode
R841 N840 N841 10
D841 N841 0 diode
R842 N841 N842 10
D842 N842 0 diode
R843 N842 N843 10
D843 N843 0 diode
R844 N843 N844 10
D844 N844 0 diode
R845 N844 N845 10
D845 N845 0 diode
R846 N845 N846 10
D846 N846 0 diode
R847 N846 N847 10
D847 N847 0 diode
R848 N847 N848 10
D848 N848 0 diode
R849 N848 N849 10
D849 N849 0 diode
R850 N849 N850 10
D850 N850 0 diode
R851 N850 N851 10
D851 N851 0 diode
R852 N851 N852 10
D852 N852 0 diode
R853 N852 N853 10
D853 N853 0 diode
R854 N853 N854 10
D854 N854 0 diode
R855 N854 N855 10
D855 N855 0 diode
R856 N855 N856 10
D856 N856 0 diode
R857 N856 N857 10
D857 N857 0 diode
R858 N857 N858 10
D858 N858 0 diode
R859 N858 N859 10
D859 N859 0 diode
R860 N859 N860 10
D860 N860 0 diode
R861 N860 N861 10
D861 N861 0 diode
R862 N861 N862 10
D862 N862 0 diode
R863 N862 N863 10
D863 N863 0 diode
R864 N863 N864 10
D864 N864 0 diode
R865 N864 N865 10
D865 N865 0 diode
R866 N865 N866 10
D866 N866 0 diode
R867 N866 N867 10
D867 N867 0 diode
R868 N867 N868 10
D868 N868 0 diode
R869 N868 N869 10
D869 N869 0 diode
R870 N869 N870 10
D870 N870 0 diode
R871 N870 N871 10
D871 N871 0 diode
R872 N871 N872 10
D872 N872 0 diode
R873 N872 N873 10
D873 N873 0 diode
R874 N873 N874 10
D874 N874 0 diode
R875 N874 N875 10
D875 N875 0 diode
R876 N875 N876 10
D876 N876 0 diode
R877 N876 N877 10
D877 N877 0 diode
R878 N877 N878 10
D878 N878 0 diode
R879 N878 N879 10
D879 N879 0 diode
R880 N879 N880 10
D880 N880 0 diode
R881 N880 N881 10
D881 N881 0 diode
R882 N881 N882 10
D882 N882 0 diode
R883 N882 N883 10
D883 N883 0 diode
R884 N883 N884 10
D884 N884 0 diode
R885 N884 N885 10
D885 N885 0 diode
R886 N885 N886 10
D886 N886 0 diode
R887 N886 N887 10
D887 N887 0 diode
R888 N887 N888 10
D888 N888 0 diode
R889 N888 N889 10
D889 N889 0 diode
R890 N889 N890 10
D890 N890 0 diode
R891 N890 N891 10
D891 N891 0 diode
R892 N891 N892 10
D892 N892 0 diode
R893 N892 N893 10
D893 N893 0 diode
R894 N893 N894 10
D894 N894 0 diode
R895 N894 N895 10
D895 N895 0 diode
R896 N895 N896 10
D896 N896 0 diode
R897 N896 N897 10
D897 N897 0 diode
R898 N897 N898 10
D898 N898 0 diode
R899 N898 N899 10
D899 N899 0 diode
R900 N899 N900 10
D900 N900 0 diode
R901 N900 N901 10
D901 N901 0 diode
R902 N901 N902 10
D902 N902 0 diode
R903 N902 N903 10
D903 N903 0 diode
R904 N903 N904 10
D904 N904 0 diode
R905 N904 N905 10
D905 N905 0 diode
R906 N905 N906 10
D906 N906 0 diode
R907 N906 N907 10
D907 N907 0 diode
R908 N907 N908 10
D908 N908 0 diode
R909 N908 N909 10
D909 N909 0 diode
R910 N909 N910 10
D910 N910 0 diode
R911 N910 N911 10
D911 N911 0 diode
R912 N911 N912 10
D912 N912 0 diode
R913 N912 N913 10
D913 N913 0 diode
R914 N913 N914 10
D914 N914 0 diode
R915 N914 N915 10
D915 N915 0 diode
R916 N915 N916 10
D916 N916 0 diode
R917 N916 N917 10
D917 N917 0 diode
R918 N917 N918 10
D918 N918 0 diode
R919 N918 N919 10
D919 N919 0 diode
R920 N919 N920 10
D920 N920 0 diode
R921 N920 N921 10
D921 N921 0 diode
R922 N921 N922 10
D922 N922 0 diode
R923 N922 N923 10
D923 N923 0 diode
R924 N923 N924 10
D924 N924 0 diode
R925 N924 N925 10
D925 N925 0 diode
R926 N925 N926 10
D926 N926 0 diode
R927 N926 N927 10
D927 N927 0 diode
R928 N927 N928 10
D928 N928 0 diode
R929 N928 N929 10
D929 N929 0 diode
R930 N929 N930 10
D930 N930 0 diode
R931 N930 N931 10
D931 N931 0 diode
R932 N931 N932 10
D932 N932 0 diode
R933 N932 N933 10
D933 N933 0 diode
R934 N933 N934 10
D934 N934 0 diode
R935 N934 N935 10
D935 N935 0 diode
R936 N935 N936 10
D936 N936 0 diode
R937 N936 N937 10
D937 N937 0 diode
R938 N937 N938 10
D938 N938 0 diode
R939 N938 N939 10
D939 N939 0 diode
R940 N939 N940 10
D940 N940 0 diode
R941 N940 N941 10
D941 N941 0 diode
R942 N941 N942 10
D942 N942 0 diode
R943 N942 N943 10
D943 N943 0 diode
R944 N943 N944 10
D944 N944 0 diode
R945 N944 N945 10
D945 N945 0 diode
R946 N945 N946 10
D946 N946 0 diode
R947 N946 N947 10
D947 N947 0 diode
R948 N947 N948 10
D948 N948 0 diode
R949 N948 N949 10
D949 N949 0 diode
R950 N949 N950 10
D950 N950 0 diode
R951 N950 N951 10
D951 N951 0 diode
R952 N951 N952 10
D952 N952 0 diode
R953 N952 N953 10
D953 N953 0 diode
R954 N953 N954 10
D954 N954 0 diode
R955 N954 N955 10
D955 N955 0 diode
R956 N955 N956 10
D956 N956 0 diode
R957 N956 N957 10
D957 N957 0 diode
R958 N957 N958 10
D958 N958 0 diode
R959 N958 N959 10
D959 N959 0 diode
R960 N959 N960 10
D960 N960 0 diode
R961 N960 N961 10
D961 N961 0 diode
R962 N961 N962 10
D962 N962 0 diode
R963 N962 N963 10
D963 N963 0 diode
R964 N963 N964 10
D964 N964 0 diode
R965 N964 N965 10
D965 N965 0 diode
R966 N965 N966 10
D966 N966 0 diode
R967 N966 N967 10
D967 N967 0 diode
R968 N967 N968 10
D968 N968 0 diode
R969 N968 N969 10
D969 N969 0 diode
R970 N969 N970 10
D970 N970 0 diode
R971 N970 N971 10
D971 N971 0 diode
R972 N971 N972 10
D972 N972 0 diode
R973 N972 N973 10
D973 N973 0 diode
R974 N973 N974 10
D974 N974 0 diode
R975 N974 N975 10
D975 N975 0 diode
R976 N975 N976 10
D976 N976 0 diode
R977 N976 N977 10
D977 N977 0 diode
R978 N977 N978 10
D978 N978 0 diode
R979 N978 N979 10
D979 N979 0 diode
R980 N979 N980 10
D980 N980 0 diode
R981 N980 N981 10
D981 N981 0 diode
R982 N981 N982 10
D982 N982 0 diode
R983 N982 N983 10
D983 N983 0 diode
R984 N983 N984 10
D984 N984 0 diode
R985 N984 N985 10
D985 N985 0 diode
R986 N985 N986 10
D986 N986 0 diode
R987 N986 N987 10
D987 N987 0 diode
R988 N987 N988 10
D988 N988 0 diode
R989 N988 N989 10
D989 N989 0 diode
R990 N989 N990 10
D990 N990 0 diode
R991 N990 N991 10
D991 N991 0 diode
R992 N991 N992 10
D992 N992 0 diode
R993 N992 N993 10
D993 N993 0 diode
R994 N993 N994 10
D994 N994 0 diode
R995 N994 N995 10
D995 N995 0 diode
R996 N995 N996 10
D996 N996 0 diode
R997 N996 N997 10
D997 N997 0 diode
R998 N997 N998 10
D998 N998 0 diode
R999 N998 N999 10
D999 N999 0 diode
R1000 N999 N1000 10
D1000 N1000 0 diode
R1001 N1000 N1001 10
D1001 N1001 0 diode
R1002 N1001 N1002 10
D1002 N1002 0 diode
R1003 N1002 N1003 10
D1003 N1003 0 diode
R1004 N1003 N1004 10
D1004 N1004 0 diode
R1005 N1004 N1005 10
D1005 N1005 0 diode
R1006 N1005 N1006 10
D1006 N1006 0 diode
R1007 N1006 N1007 10
D1007 N1007 0 diode
R1008 N1007 N1008 10
D1008 N1008 0 diode
R1009 N1008 N1009 10
D1009 N1009 0 diode
R1010 N1009 N1010 10
D1010 N1010 0 diode
R1011 N1010 N1011 10
D1011 N1011 0 diode
R1012 N1011 N1012 10
D1012 N1012 0 diode
R1013 N1012 N1013 10
D1013 N1013 0 diode
R1014 N1013 N1014 10
D1014 N1014 0 diode
R1015 N1014 N1015 10
D1015 N1015 0 diode
R1016 N1015 N1016 10
D1016 N1016 0 diode
R1017 N1016 N1017 10
D1017 N1017 0 diode
R1018 N1017 N1018 10
D1018 N1018 0 diode
R1019 N1018 N1019 10
D1019 N1019 0 diode
R1020 N1019 N1020 10
D1020 N1020 0 diode
R1021 N1020 N1021 10
D1021 N1021 0 diode
R1022 N1021 N1022 10
D1022 N1022 0 diode
R1023 N1022 N1023 10
D1023 N1023 0 diode
R1024 N1023 N1024 10
D1024 N1024 0 diode
R1025 N1024 N1025 10
D1025 N1025 0 diode
R1026 N1025 N1026 10
D1026 N1026 0 diode
R1027 N1026 N1027 10
D1027 N1027 0 diode
R1028 N1027 N1028 10
D1028 N1028 0 diode
R1029 N1028 N1029 10
D1029 N1029 0 diode
R1030 N1029 N1030 10
D1030 N1030 0 diode
R1031 N1030 N1031 10
D1031 N1031 0 diode
R1032 N1031 N1032 10
D1032 N1032 0 diode
R1033 N1032 N1033 10
D1033 N1033 0 diode
R1034 N1033 N1034 10
D1034 N1034 0 diode
R1035 N1034 N1035 10
D1035 N1035 0 diode
R1036 N1035 N1036 10
D1036 N1036 0 diode
R1037 N1036 N1037 10
D1037 N1037 0 diode
R1038 N1037 N1038 10
D1038 N1038 0 diode
R1039 N1038 N1039 10
D1039 N1039 0 diode
R1040 N1039 N1040 10
D1040 N1040 0 diode
R1041 N1040 N1041 10
D1041 N1041 0 diode
R1042 N1041 N1042 10
D1042 N1042 0 diode
R1043 N1042 N1043 10
D1043 N1043 0 diode
R1044 N1043 N1044 10
D1044 N1044 0 diode
R1045 N1044 N1045 10
D1045 N1045 0 diode
R1046 N1045 N1046 10
D1046 N1046 0 diode
R1047 N1046 N1047 10
D1047 N1047 0 diode
R1048 N1047 N1048 10
D1048 N1048 0 diode
R1049 N1048 N1049 10
D1049 N1049 0 diode
R1050 N1049 N1050 10
D1050 N1050 0 diode
R1051 N1050 N1051 10
D1051 N1051 0 diode
R1052 N1051 N1052 10
D1052 N1052 0 diode
R1053 N1052 N1053 10
D1053 N1053 0 diode
R1054 N1053 N1054 10
D1054 N1054 0 diode
R1055 N1054 N1055 10
D1055 N1055 0 diode
R1056 N1055 N1056 10
D1056 N1056 0 diode
R1057 N1056 N1057 10
D1057 N1057 0 diode
R1058 N1057 N1058 10
D1058 N1058 0 diode
R1059 N1058 N1059 10
D1059 N1059 0 diode
R1060 N1059 N1060 10
D1060 N1060 0 diode
R1061 N1060 N1061 10
D1061 N1061 0 diode
R1062 N1061 N1062 10
D1062 N1062 0 diode
R1063 N1062 N1063 10
D1063 N1063 0 diode
R1064 N1063 N1064 10
D1064 N1064 0 diode
R1065 N1064 N1065 10
D1065 N1065 0 diode
R1066 N1065 N1066 10
D1066 N1066 0 diode
R1067 N1066 N1067 10
D1067 N1067 0 diode
R1068 N1067 N1068 10
D1068 N1068 0 diode
R1069 N1068 N1069 10
D1069 N1069 0 diode
R1070 N1069 N1070 10
D1070 N1070 0 diode
R1071 N1070 N1071 10
D1071 N1071 0 diode
R1072 N1071 N1072 10
D1072 N1072 0 diode
R1073 N1072 N1073 10
D1073 N1073 0 diode
R1074 N1073 N1074 10
D1074 N1074 0 diode
R1075 N1074 N1075 10
D1075 N1075 0 diode
R1076 N1075 N1076 10
D1076 N1076 0 diode
R1077 N1076 N1077 10
D1077 N1077 0 diode
R1078 N1077 N1078 10
D1078 N1078 0 diode
R1079 N1078 N1079 10
D1079 N1079 0 diode
R1080 N1079 N1080 10
D1080 N1080 0 diode
R1081 N1080 N1081 10
D1081 N1081 0 diode
R1082 N1081 N1082 10
D1082 N1082 0 diode
R1083 N1082 N1083 10
D1083 N1083 0 diode
R1084 N1083 N1084 10
D1084 N1084 0 diode
R1085 N1084 N1085 10
D1085 N1085 0 diode
R1086 N1085 N1086 10
D1086 N1086 0 diode
R1087 N1086 N1087 10
D1087 N1087 0 diode
R1088 N1087 N1088 10
D1088 N1088 0 diode
R1089 N1088 N1089 10
D1089 N1089 0 diode
R1090 N1089 N1090 10
D1090 N1090 0 diode
R1091 N1090 N1091 10
D1091 N1091 0 diode
R1092 N1091 N1092 10
D1092 N1092 0 diode
R1093 N1092 N1093 10
D1093 N1093 0 diode
R1094 N1093 N1094 10
D1094 N1094 0 diode
R1095 N1094 N1095 10
D1095 N1095 0 diode
R1096 N1095 N1096 10
D1096 N1096 0 diode
R1097 N1096 N1097 10
D1097 N1097 0 diode
R1098 N1097 N1098 10
D1098 N1098 0 diode
R1099 N1098 N1099 10
D1099 N1099 0 diode
R1100 N1099 N1100 10
D1100 N1100 0 diode
R1101 N1100 N1101 10
D1101 N1101 0 diode
R1102 N1101 N1102 10
D1102 N1102 0 diode
R1103 N1102 N1103 10
D1103 N1103 0 diode
R1104 N1103 N1104 10
D1104 N1104 0 diode
R1105 N1104 N1105 10
D1105 N1105 0 diode
R1106 N1105 N1106 10
D1106 N1106 0 diode
R1107 N1106 N1107 10
D1107 N1107 0 diode
R1108 N1107 N1108 10
D1108 N1108 0 diode
R1109 N1108 N1109 10
D1109 N1109 0 diode
R1110 N1109 N1110 10
D1110 N1110 0 diode
R1111 N1110 N1111 10
D1111 N1111 0 diode
R1112 N1111 N1112 10
D1112 N1112 0 diode
R1113 N1112 N1113 10
D1113 N1113 0 diode
R1114 N1113 N1114 10
D1114 N1114 0 diode
R1115 N1114 N1115 10
D1115 N1115 0 diode
R1116 N1115 N1116 10
D1116 N1116 0 diode
R1117 N1116 N1117 10
D1117 N1117 0 diode
R1118 N1117 N1118 10
D1118 N1118 0 diode
R1119 N1118 N1119 10
D1119 N1119 0 diode
R1120 N1119 N1120 10
D1120 N1120 0 diode
R1121 N1120 N1121 10
D1121 N1121 0 diode
R1122 N1121 N1122 10
D1122 N1122 0 diode
R1123 N1122 N1123 10
D1123 N1123 0 diode
R1124 N1123 N1124 10
D1124 N1124 0 diode
R1125 N1124 N1125 10
D1125 N1125 0 diode
R1126 N1125 N1126 10
D1126 N1126 0 diode
R1127 N1126 N1127 10
D1127 N1127 0 diode
R1128 N1127 N1128 10
D1128 N1128 0 diode
R1129 N1128 N1129 10
D1129 N1129 0 diode
R1130 N1129 N1130 10
D1130 N1130 0 diode
R1131 N1130 N1131 10
D1131 N1131 0 diode
R1132 N1131 N1132 10
D1132 N1132 0 diode
R1133 N1132 N1133 10
D1133 N1133 0 diode
R1134 N1133 N1134 10
D1134 N1134 0 diode
R1135 N1134 N1135 10
D1135 N1135 0 diode
R1136 N1135 N1136 10
D1136 N1136 0 diode
R1137 N1136 N1137 10
D1137 N1137 0 diode
R1138 N1137 N1138 10
D1138 N1138 0 diode
R1139 N1138 N1139 10
D1139 N1139 0 diode
R1140 N1139 N1140 10
D1140 N1140 0 diode
R1141 N1140 N1141 10
D1141 N1141 0 diode
R1142 N1141 N1142 10
D1142 N1142 0 diode
R1143 N1142 N1143 10
D1143 N1143 0 diode
R1144 N1143 N1144 10
D1144 N1144 0 diode
R1145 N1144 N1145 10
D1145 N1145 0 diode
R1146 N1145 N1146 10
D1146 N1146 0 diode
R1147 N1146 N1147 10
D1147 N1147 0 diode
R1148 N1147 N1148 10
D1148 N1148 0 diode
R1149 N1148 N1149 10
D1149 N1149 0 diode
R1150 N1149 N1150 10
D1150 N1150 0 diode
R1151 N1150 N1151 10
D1151 N1151 0 diode
R1152 N1151 N1152 10
D1152 N1152 0 diode
R1153 N1152 N1153 10
D1153 N1153 0 diode
R1154 N1153 N1154 10
D1154 N1154 0 diode
R1155 N1154 N1155 10
D1155 N1155 0 diode
R1156 N1155 N1156 10
D1156 N1156 0 diode
R1157 N1156 N1157 10
D1157 N1157 0 diode
R1158 N1157 N1158 10
D1158 N1158 0 diode
R1159 N1158 N1159 10
D1159 N1159 0 diode
R1160 N1159 N1160 10
D1160 N1160 0 diode
R1161 N1160 N1161 10
D1161 N1161 0 diode
R1162 N1161 N1162 10
D1162 N1162 0 diode
R1163 N1162 N1163 10
D1163 N1163 0 diode
R1164 N1163 N1164 10
D1164 N1164 0 diode
R1165 N1164 N1165 10
D1165 N1165 0 diode
R1166 N1165 N1166 10
D1166 N1166 0 diode
R1167 N1166 N1167 10
D1167 N1167 0 diode
R1168 N1167 N1168 10
D1168 N1168 0 diode
R1169 N1168 N1169 10
D1169 N1169 0 diode
R1170 N1169 N1170 10
D1170 N1170 0 diode
R1171 N1170 N1171 10
D1171 N1171 0 diode
R1172 N1171 N1172 10
D1172 N1172 0 diode
R1173 N1172 N1173 10
D1173 N1173 0 diode
R1174 N1173 N1174 10
D1174 N1174 0 diode
R1175 N1174 N1175 10
D1175 N1175 0 diode
R1176 N1175 N1176 10
D1176 N1176 0 diode
R1177 N1176 N1177 10
D1177 N1177 0 diode
R1178 N1177 N1178 10
D1178 N1178 0 diode
R1179 N1178 N1179 10
D1179 N1179 0 diode
R1180 N1179 N1180 10
D1180 N1180 0 diode
R1181 N1180 N1181 10
D1181 N1181 0 diode
R1182 N1181 N1182 10
D1182 N1182 0 diode
R1183 N1182 N1183 10
D1183 N1183 0 diode
R1184 N1183 N1184 10
D1184 N1184 0 diode
R1185 N1184 N1185 10
D1185 N1185 0 diode
R1186 N1185 N1186 10
D1186 N1186 0 diode
R1187 N1186 N1187 10
D1187 N1187 0 diode
R1188 N1187 N1188 10
D1188 N1188 0 diode
R1189 N1188 N1189 10
D1189 N1189 0 diode
R1190 N1189 N1190 10
D1190 N1190 0 diode
R1191 N1190 N1191 10
D1191 N1191 0 diode
R1192 N1191 N1192 10
D1192 N1192 0 diode
R1193 N1192 N1193 10
D1193 N1193 0 diode
R1194 N1193 N1194 10
D1194 N1194 0 diode
R1195 N1194 N1195 10
D1195 N1195 0 diode
R1196 N1195 N1196 10
D1196 N1196 0 diode
R1197 N1196 N1197 10
D1197 N1197 0 diode
R1198 N1197 N1198 10
D1198 N1198 0 diode
R1199 N1198 N1199 10
D1199 N1199 0 diode
R1200 N1199 N1200 10
D1200 N1200 0 diode
R1201 N1200 N1201 10
D1201 N1201 0 diode
R1202 N1201 N1202 10
D1202 N1202 0 diode
R1203 N1202 N1203 10
D1203 N1203 0 diode
R1204 N1203 N1204 10
D1204 N1204 0 diode
R1205 N1204 N1205 10
D1205 N1205 0 diode
R1206 N1205 N1206 10
D1206 N1206 0 diode
R1207 N1206 N1207 10
D1207 N1207 0 diode
R1208 N1207 N1208 10
D1208 N1208 0 diode
R1209 N1208 N1209 10
D1209 N1209 0 diode
R1210 N1209 N1210 10
D1210 N1210 0 diode
R1211 N1210 N1211 10
D1211 N1211 0 diode
R1212 N1211 N1212 10
D1212 N1212 0 diode
R1213 N1212 N1213 10
D1213 N1213 0 diode
R1214 N1213 N1214 10
D1214 N1214 0 diode
R1215 N1214 N1215 10
D1215 N1215 0 diode
R1216 N1215 N1216 10
D1216 N1216 0 diode
R1217 N1216 N1217 10
D1217 N1217 0 diode
R1218 N1217 N1218 10
D1218 N1218 0 diode
R1219 N1218 N1219 10
D1219 N1219 0 diode
R1220 N1219 N1220 10
D1220 N1220 0 diode
R1221 N1220 N1221 10
D1221 N1221 0 diode
R1222 N1221 N1222 10
D1222 N1222 0 diode
R1223 N1222 N1223 10
D1223 N1223 0 diode
R1224 N1223 N1224 10
D1224 N1224 0 diode
R1225 N1224 N1225 10
D1225 N1225 0 diode
R1226 N1225 N1226 10
D1226 N1226 0 diode
R1227 N1226 N1227 10
D1227 N1227 0 diode
R1228 N1227 N1228 10
D1228 N1228 0 diode
R1229 N1228 N1229 10
D1229 N1229 0 diode
R1230 N1229 N1230 10
D1230 N1230 0 diode
R1231 N1230 N1231 10
D1231 N1231 0 diode
R1232 N1231 N1232 10
D1232 N1232 0 diode
R1233 N1232 N1233 10
D1233 N1233 0 diode
R1234 N1233 N1234 10
D1234 N1234 0 diode
R1235 N1234 N1235 10
D1235 N1235 0 diode
R1236 N1235 N1236 10
D1236 N1236 0 diode
R1237 N1236 N1237 10
D1237 N1237 0 diode
R1238 N1237 N1238 10
D1238 N1238 0 diode
R1239 N1238 N1239 10
D1239 N1239 0 diode
R1240 N1239 N1240 10
D1240 N1240 0 diode
R1241 N1240 N1241 10
D1241 N1241 0 diode
R1242 N1241 N1242 10
D1242 N1242 0 diode
R1243 N1242 N1243 10
D1243 N1243 0 diode
R1244 N1243 N1244 10
D1244 N1244 0 diode
R1245 N1244 N1245 10
D1245 N1245 0 diode
R1246 N1245 N1246 10
D1246 N1246 0 diode
R1247 N1246 N1247 10
D1247 N1247 0 diode
R1248 N1247 N1248 10
D1248 N1248 0 diode
R1249 N1248 N1249 10
D1249 N1249 0 diode
R1250 N1249 N1250 10
D1250 N1250 0 diode
R1251 N1250 N1251 10
D1251 N1251 0 diode
R1252 N1251 N1252 10
D1252 N1252 0 diode
R1253 N1252 N1253 10
D1253 N1253 0 diode
R1254 N1253 N1254 10
D1254 N1254 0 diode
R1255 N1254 N1255 10
D1255 N1255 0 diode
R1256 N1255 N1256 10
D1256 N1256 0 diode
R1257 N1256 N1257 10
D1257 N1257 0 diode
R1258 N1257 N1258 10
D1258 N1258 0 diode
R1259 N1258 N1259 10
D1259 N1259 0 diode
R1260 N1259 N1260 10
D1260 N1260 0 diode
R1261 N1260 N1261 10
D1261 N1261 0 diode
R1262 N1261 N1262 10
D1262 N1262 0 diode
R1263 N1262 N1263 10
D1263 N1263 0 diode
R1264 N1263 N1264 10
D1264 N1264 0 diode
R1265 N1264 N1265 10
D1265 N1265 0 diode
R1266 N1265 N1266 10
D1266 N1266 0 diode
R1267 N1266 N1267 10
D1267 N1267 0 diode
R1268 N1267 N1268 10
D1268 N1268 0 diode
R1269 N1268 N1269 10
D1269 N1269 0 diode
R1270 N1269 N1270 10
D1270 N1270 0 diode
R1271 N1270 N1271 10
D1271 N1271 0 diode
R1272 N1271 N1272 10
D1272 N1272 0 diode
R1273 N1272 N1273 10
D1273 N1273 0 diode
R1274 N1273 N1274 10
D1274 N1274 0 diode
R1275 N1274 N1275 10
D1275 N1275 0 diode
R1276 N1275 N1276 10
D1276 N1276 0 diode
R1277 N1276 N1277 10
D1277 N1277 0 diode
R1278 N1277 N1278 10
D1278 N1278 0 diode
R1279 N1278 N1279 10
D1279 N1279 0 diode
R1280 N1279 N1280 10
D1280 N1280 0 diode
R1281 N1280 N1281 10
D1281 N1281 0 diode
R1282 N1281 N1282 10
D1282 N1282 0 diode
R1283 N1282 N1283 10
D1283 N1283 0 diode
R1284 N1283 N1284 10
D1284 N1284 0 diode
R1285 N1284 N1285 10
D1285 N1285 0 diode
R1286 N1285 N1286 10
D1286 N1286 0 diode
R1287 N1286 N1287 10
D1287 N1287 0 diode
R1288 N1287 N1288 10
D1288 N1288 0 diode
R1289 N1288 N1289 10
D1289 N1289 0 diode
R1290 N1289 N1290 10
D1290 N1290 0 diode
R1291 N1290 N1291 10
D1291 N1291 0 diode
R1292 N1291 N1292 10
D1292 N1292 0 diode
R1293 N1292 N1293 10
D1293 N1293 0 diode
R1294 N1293 N1294 10
D1294 N1294 0 diode
R1295 N1294 N1295 10
D1295 N1295 0 diode
R1296 N1295 N1296 10
D1296 N1296 0 diode
R1297 N1296 N1297 10
D1297 N1297 0 diode
R1298 N1297 N1298 10
D1298 N1298 0 diode
R1299 N1298 N1299 10
D1299 N1299 0 diode
R1300 N1299 N1300 10
D1300 N1300 0 diode
R1301 N1300 N1301 10
D1301 N1301 0 diode
R1302 N1301 N1302 10
D1302 N1302 0 diode
R1303 N1302 N1303 10
D1303 N1303 0 diode
R1304 N1303 N1304 10
D1304 N1304 0 diode
R1305 N1304 N1305 10
D1305 N1305 0 diode
R1306 N1305 N1306 10
D1306 N1306 0 diode
R1307 N1306 N1307 10
D1307 N1307 0 diode
R1308 N1307 N1308 10
D1308 N1308 0 diode
R1309 N1308 N1309 10
D1309 N1309 0 diode
R1310 N1309 N1310 10
D1310 N1310 0 diode
R1311 N1310 N1311 10
D1311 N1311 0 diode
R1312 N1311 N1312 10
D1312 N1312 0 diode
R1313 N1312 N1313 10
D1313 N1313 0 diode
R1314 N1313 N1314 10
D1314 N1314 0 diode
R1315 N1314 N1315 10
D1315 N1315 0 diode
R1316 N1315 N1316 10
D1316 N1316 0 diode
R1317 N1316 N1317 10
D1317 N1317 0 diode
R1318 N1317 N1318 10
D1318 N1318 0 diode
R1319 N1318 N1319 10
D1319 N1319 0 diode
R1320 N1319 N1320 10
D1320 N1320 0 diode
R1321 N1320 N1321 10
D1321 N1321 0 diode
R1322 N1321 N1322 10
D1322 N1322 0 diode
R1323 N1322 N1323 10
D1323 N1323 0 diode
R1324 N1323 N1324 10
D1324 N1324 0 diode
R1325 N1324 N1325 10
D1325 N1325 0 diode
R1326 N1325 N1326 10
D1326 N1326 0 diode
R1327 N1326 N1327 10
D1327 N1327 0 diode
R1328 N1327 N1328 10
D1328 N1328 0 diode
R1329 N1328 N1329 10
D1329 N1329 0 diode
R1330 N1329 N1330 10
D1330 N1330 0 diode
R1331 N1330 N1331 10
D1331 N1331 0 diode
R1332 N1331 N1332 10
D1332 N1332 0 diode
R1333 N1332 N1333 10
D1333 N1333 0 diode
R1334 N1333 N1334 10
D1334 N1334 0 diode
R1335 N1334 N1335 10
D1335 N1335 0 diode
R1336 N1335 N1336 10
D1336 N1336 0 diode
R1337 N1336 N1337 10
D1337 N1337 0 diode
R1338 N1337 N1338 10
D1338 N1338 0 diode
R1339 N1338 N1339 10
D1339 N1339 0 diode
R1340 N1339 N1340 10
D1340 N1340 0 diode
R1341 N1340 N1341 10
D1341 N1341 0 diode
R1342 N1341 N1342 10
D1342 N1342 0 diode
R1343 N1342 N1343 10
D1343 N1343 0 diode
R1344 N1343 N1344 10
D1344 N1344 0 diode
R1345 N1344 N1345 10
D1345 N1345 0 diode
R1346 N1345 N1346 10
D1346 N1346 0 diode
R1347 N1346 N1347 10
D1347 N1347 0 diode
R1348 N1347 N1348 10
D1348 N1348 0 diode
R1349 N1348 N1349 10
D1349 N1349 0 diode
R1350 N1349 N1350 10
D1350 N1350 0 diode
R1351 N1350 N1351 10
D1351 N1351 0 diode
R1352 N1351 N1352 10
D1352 N1352 0 diode
R1353 N1352 N1353 10
D1353 N1353 0 diode
R1354 N1353 N1354 10
D1354 N1354 0 diode
R1355 N1354 N1355 10
D1355 N1355 0 diode
R1356 N1355 N1356 10
D1356 N1356 0 diode
R1357 N1356 N1357 10
D1357 N1357 0 diode
R1358 N1357 N1358 10
D1358 N1358 0 diode
R1359 N1358 N1359 10
D1359 N1359 0 diode
R1360 N1359 N1360 10
D1360 N1360 0 diode
R1361 N1360 N1361 10
D1361 N1361 0 diode
R1362 N1361 N1362 10
D1362 N1362 0 diode
R1363 N1362 N1363 10
D1363 N1363 0 diode
R1364 N1363 N1364 10
D1364 N1364 0 diode
R1365 N1364 N1365 10
D1365 N1365 0 diode
R1366 N1365 N1366 10
D1366 N1366 0 diode
R1367 N1366 N1367 10
D1367 N1367 0 diode
R1368 N1367 N1368 10
D1368 N1368 0 diode
R1369 N1368 N1369 10
D1369 N1369 0 diode
R1370 N1369 N1370 10
D1370 N1370 0 diode
R1371 N1370 N1371 10
D1371 N1371 0 diode
R1372 N1371 N1372 10
D1372 N1372 0 diode
R1373 N1372 N1373 10
D1373 N1373 0 diode
R1374 N1373 N1374 10
D1374 N1374 0 diode
R1375 N1374 N1375 10
D1375 N1375 0 diode
R1376 N1375 N1376 10
D1376 N1376 0 diode
R1377 N1376 N1377 10
D1377 N1377 0 diode
R1378 N1377 N1378 10
D1378 N1378 0 diode
R1379 N1378 N1379 10
D1379 N1379 0 diode
R1380 N1379 N1380 10
D1380 N1380 0 diode
R1381 N1380 N1381 10
D1381 N1381 0 diode
R1382 N1381 N1382 10
D1382 N1382 0 diode
R1383 N1382 N1383 10
D1383 N1383 0 diode
R1384 N1383 N1384 10
D1384 N1384 0 diode
R1385 N1384 N1385 10
D1385 N1385 0 diode
R1386 N1385 N1386 10
D1386 N1386 0 diode
R1387 N1386 N1387 10
D1387 N1387 0 diode
R1388 N1387 N1388 10
D1388 N1388 0 diode
R1389 N1388 N1389 10
D1389 N1389 0 diode
R1390 N1389 N1390 10
D1390 N1390 0 diode
R1391 N1390 N1391 10
D1391 N1391 0 diode
R1392 N1391 N1392 10
D1392 N1392 0 diode
R1393 N1392 N1393 10
D1393 N1393 0 diode
R1394 N1393 N1394 10
D1394 N1394 0 diode
R1395 N1394 N1395 10
D1395 N1395 0 diode
R1396 N1395 N1396 10
D1396 N1396 0 diode
R1397 N1396 N1397 10
D1397 N1397 0 diode
R1398 N1397 N1398 10
D1398 N1398 0 diode
R1399 N1398 N1399 10
D1399 N1399 0 diode
R1400 N1399 N1400 10
D1400 N1400 0 diode
R1401 N1400 N1401 10
D1401 N1401 0 diode
R1402 N1401 N1402 10
D1402 N1402 0 diode
R1403 N1402 N1403 10
D1403 N1403 0 diode
R1404 N1403 N1404 10
D1404 N1404 0 diode
R1405 N1404 N1405 10
D1405 N1405 0 diode
R1406 N1405 N1406 10
D1406 N1406 0 diode
R1407 N1406 N1407 10
D1407 N1407 0 diode
R1408 N1407 N1408 10
D1408 N1408 0 diode
R1409 N1408 N1409 10
D1409 N1409 0 diode
R1410 N1409 N1410 10
D1410 N1410 0 diode
R1411 N1410 N1411 10
D1411 N1411 0 diode
R1412 N1411 N1412 10
D1412 N1412 0 diode
R1413 N1412 N1413 10
D1413 N1413 0 diode
R1414 N1413 N1414 10
D1414 N1414 0 diode
R1415 N1414 N1415 10
D1415 N1415 0 diode
R1416 N1415 N1416 10
D1416 N1416 0 diode
R1417 N1416 N1417 10
D1417 N1417 0 diode
R1418 N1417 N1418 10
D1418 N1418 0 diode
R1419 N1418 N1419 10
D1419 N1419 0 diode
R1420 N1419 N1420 10
D1420 N1420 0 diode
R1421 N1420 N1421 10
D1421 N1421 0 diode
R1422 N1421 N1422 10
D1422 N1422 0 diode
R1423 N1422 N1423 10
D1423 N1423 0 diode
R1424 N1423 N1424 10
D1424 N1424 0 diode
R1425 N1424 N1425 10
D1425 N1425 0 diode
R1426 N1425 N1426 10
D1426 N1426 0 diode
R1427 N1426 N1427 10
D1427 N1427 0 diode
R1428 N1427 N1428 10
D1428 N1428 0 diode
R1429 N1428 N1429 10
D1429 N1429 0 diode
R1430 N1429 N1430 10
D1430 N1430 0 diode
R1431 N1430 N1431 10
D1431 N1431 0 diode
R1432 N1431 N1432 10
D1432 N1432 0 diode
R1433 N1432 N1433 10
D1433 N1433 0 diode
R1434 N1433 N1434 10
D1434 N1434 0 diode
R1435 N1434 N1435 10
D1435 N1435 0 diode
R1436 N1435 N1436 10
D1436 N1436 0 diode
R1437 N1436 N1437 10
D1437 N1437 0 diode
R1438 N1437 N1438 10
D1438 N1438 0 diode
R1439 N1438 N1439 10
D1439 N1439 0 diode
R1440 N1439 N1440 10
D1440 N1440 0 diode
R1441 N1440 N1441 10
D1441 N1441 0 diode
R1442 N1441 N1442 10
D1442 N1442 0 diode
R1443 N1442 N1443 10
D1443 N1443 0 diode
R1444 N1443 N1444 10
D1444 N1444 0 diode
R1445 N1444 N1445 10
D1445 N1445 0 diode
R1446 N1445 N1446 10
D1446 N1446 0 diode
R1447 N1446 N1447 10
D1447 N1447 0 diode
R1448 N1447 N1448 10
D1448 N1448 0 diode
R1449 N1448 N1449 10
D1449 N1449 0 diode
R1450 N1449 N1450 10
D1450 N1450 0 diode
R1451 N1450 N1451 10
D1451 N1451 0 diode
R1452 N1451 N1452 10
D1452 N1452 0 diode
R1453 N1452 N1453 10
D1453 N1453 0 diode
R1454 N1453 N1454 10
D1454 N1454 0 diode
R1455 N1454 N1455 10
D1455 N1455 0 diode
R1456 N1455 N1456 10
D1456 N1456 0 diode
R1457 N1456 N1457 10
D1457 N1457 0 diode
R1458 N1457 N1458 10
D1458 N1458 0 diode
R1459 N1458 N1459 10
D1459 N1459 0 diode
R1460 N1459 N1460 10
D1460 N1460 0 diode
R1461 N1460 N1461 10
D1461 N1461 0 diode
R1462 N1461 N1462 10
D1462 N1462 0 diode
R1463 N1462 N1463 10
D1463 N1463 0 diode
R1464 N1463 N1464 10
D1464 N1464 0 diode
R1465 N1464 N1465 10
D1465 N1465 0 diode
R1466 N1465 N1466 10
D1466 N1466 0 diode
R1467 N1466 N1467 10
D1467 N1467 0 diode
R1468 N1467 N1468 10
D1468 N1468 0 diode
R1469 N1468 N1469 10
D1469 N1469 0 diode
R1470 N1469 N1470 10
D1470 N1470 0 diode
R1471 N1470 N1471 10
D1471 N1471 0 diode
R1472 N1471 N1472 10
D1472 N1472 0 diode
R1473 N1472 N1473 10
D1473 N1473 0 diode
R1474 N1473 N1474 10
D1474 N1474 0 diode
R1475 N1474 N1475 10
D1475 N1475 0 diode
R1476 N1475 N1476 10
D1476 N1476 0 diode
R1477 N1476 N1477 10
D1477 N1477 0 diode
R1478 N1477 N1478 10
D1478 N1478 0 diode
R1479 N1478 N1479 10
D1479 N1479 0 diode
R1480 N1479 N1480 10
D1480 N1480 0 diode
R1481 N1480 N1481 10
D1481 N1481 0 diode
R1482 N1481 N1482 10
D1482 N1482 0 diode
R1483 N1482 N1483 10
D1483 N1483 0 diode
R1484 N1483 N1484 10
D1484 N1484 0 diode
R1485 N1484 N1485 10
D1485 N1485 0 diode
R1486 N1485 N1486 10
D1486 N1486 0 diode
R1487 N1486 N1487 10
D1487 N1487 0 diode
R1488 N1487 N1488 10
D1488 N1488 0 diode
R1489 N1488 N1489 10
D1489 N1489 0 diode
R1490 N1489 N1490 10
D1490 N1490 0 diode
R1491 N1490 N1491 10
D1491 N1491 0 diode
R1492 N1491 N1492 10
D1492 N1492 0 diode
R1493 N1492 N1493 10
D1493 N1493 0 diode
R1494 N1493 N1494 10
D1494 N1494 0 diode
R1495 N1494 N1495 10
D1495 N1495 0 diode
R1496 N1495 N1496 10
D1496 N1496 0 diode
R1497 N1496 N1497 10
D1497 N1497 0 diode
R1498 N1497 N1498 10
D1498 N1498 0 diode
R1499 N1498 N1499 10
D1499 N1499 0 diode
R1500 N1499 N1500 10
D1500 N1500 0 diode
R1501 N1500 N1501 10
D1501 N1501 0 diode
R1502 N1501 N1502 10
D1502 N1502 0 diode
R1503 N1502 N1503 10
D1503 N1503 0 diode
R1504 N1503 N1504 10
D1504 N1504 0 diode
R1505 N1504 N1505 10
D1505 N1505 0 diode
R1506 N1505 N1506 10
D1506 N1506 0 diode
R1507 N1506 N1507 10
D1507 N1507 0 diode
R1508 N1507 N1508 10
D1508 N1508 0 diode
R1509 N1508 N1509 10
D1509 N1509 0 diode
R1510 N1509 N1510 10
D1510 N1510 0 diode
R1511 N1510 N1511 10
D1511 N1511 0 diode
R1512 N1511 N1512 10
D1512 N1512 0 diode
R1513 N1512 N1513 10
D1513 N1513 0 diode
R1514 N1513 N1514 10
D1514 N1514 0 diode
R1515 N1514 N1515 10
D1515 N1515 0 diode
R1516 N1515 N1516 10
D1516 N1516 0 diode
R1517 N1516 N1517 10
D1517 N1517 0 diode
R1518 N1517 N1518 10
D1518 N1518 0 diode
R1519 N1518 N1519 10
D1519 N1519 0 diode
R1520 N1519 N1520 10
D1520 N1520 0 diode
R1521 N1520 N1521 10
D1521 N1521 0 diode
R1522 N1521 N1522 10
D1522 N1522 0 diode
R1523 N1522 N1523 10
D1523 N1523 0 diode
R1524 N1523 N1524 10
D1524 N1524 0 diode
R1525 N1524 N1525 10
D1525 N1525 0 diode
R1526 N1525 N1526 10
D1526 N1526 0 diode
R1527 N1526 N1527 10
D1527 N1527 0 diode
R1528 N1527 N1528 10
D1528 N1528 0 diode
R1529 N1528 N1529 10
D1529 N1529 0 diode
R1530 N1529 N1530 10
D1530 N1530 0 diode
R1531 N1530 N1531 10
D1531 N1531 0 diode
R1532 N1531 N1532 10
D1532 N1532 0 diode
R1533 N1532 N1533 10
D1533 N1533 0 diode
R1534 N1533 N1534 10
D1534 N1534 0 diode
R1535 N1534 N1535 10
D1535 N1535 0 diode
R1536 N1535 N1536 10
D1536 N1536 0 diode
R1537 N1536 N1537 10
D1537 N1537 0 diode
R1538 N1537 N1538 10
D1538 N1538 0 diode
R1539 N1538 N1539 10
D1539 N1539 0 diode
R1540 N1539 N1540 10
D1540 N1540 0 diode
R1541 N1540 N1541 10
D1541 N1541 0 diode
R1542 N1541 N1542 10
D1542 N1542 0 diode
R1543 N1542 N1543 10
D1543 N1543 0 diode
R1544 N1543 N1544 10
D1544 N1544 0 diode
R1545 N1544 N1545 10
D1545 N1545 0 diode
R1546 N1545 N1546 10
D1546 N1546 0 diode
R1547 N1546 N1547 10
D1547 N1547 0 diode
R1548 N1547 N1548 10
D1548 N1548 0 diode
R1549 N1548 N1549 10
D1549 N1549 0 diode
R1550 N1549 N1550 10
D1550 N1550 0 diode
R1551 N1550 N1551 10
D1551 N1551 0 diode
R1552 N1551 N1552 10
D1552 N1552 0 diode
R1553 N1552 N1553 10
D1553 N1553 0 diode
R1554 N1553 N1554 10
D1554 N1554 0 diode
R1555 N1554 N1555 10
D1555 N1555 0 diode
R1556 N1555 N1556 10
D1556 N1556 0 diode
R1557 N1556 N1557 10
D1557 N1557 0 diode
R1558 N1557 N1558 10
D1558 N1558 0 diode
R1559 N1558 N1559 10
D1559 N1559 0 diode
R1560 N1559 N1560 10
D1560 N1560 0 diode
R1561 N1560 N1561 10
D1561 N1561 0 diode
R1562 N1561 N1562 10
D1562 N1562 0 diode
R1563 N1562 N1563 10
D1563 N1563 0 diode
R1564 N1563 N1564 10
D1564 N1564 0 diode
R1565 N1564 N1565 10
D1565 N1565 0 diode
R1566 N1565 N1566 10
D1566 N1566 0 diode
R1567 N1566 N1567 10
D1567 N1567 0 diode
R1568 N1567 N1568 10
D1568 N1568 0 diode
R1569 N1568 N1569 10
D1569 N1569 0 diode
R1570 N1569 N1570 10
D1570 N1570 0 diode
R1571 N1570 N1571 10
D1571 N1571 0 diode
R1572 N1571 N1572 10
D1572 N1572 0 diode
R1573 N1572 N1573 10
D1573 N1573 0 diode
R1574 N1573 N1574 10
D1574 N1574 0 diode
R1575 N1574 N1575 10
D1575 N1575 0 diode
R1576 N1575 N1576 10
D1576 N1576 0 diode
R1577 N1576 N1577 10
D1577 N1577 0 diode
R1578 N1577 N1578 10
D1578 N1578 0 diode
R1579 N1578 N1579 10
D1579 N1579 0 diode
R1580 N1579 N1580 10
D1580 N1580 0 diode
R1581 N1580 N1581 10
D1581 N1581 0 diode
R1582 N1581 N1582 10
D1582 N1582 0 diode
R1583 N1582 N1583 10
D1583 N1583 0 diode
R1584 N1583 N1584 10
D1584 N1584 0 diode
R1585 N1584 N1585 10
D1585 N1585 0 diode
R1586 N1585 N1586 10
D1586 N1586 0 diode
R1587 N1586 N1587 10
D1587 N1587 0 diode
R1588 N1587 N1588 10
D1588 N1588 0 diode
R1589 N1588 N1589 10
D1589 N1589 0 diode
R1590 N1589 N1590 10
D1590 N1590 0 diode
R1591 N1590 N1591 10
D1591 N1591 0 diode
R1592 N1591 N1592 10
D1592 N1592 0 diode
R1593 N1592 N1593 10
D1593 N1593 0 diode
R1594 N1593 N1594 10
D1594 N1594 0 diode
R1595 N1594 N1595 10
D1595 N1595 0 diode
R1596 N1595 N1596 10
D1596 N1596 0 diode
R1597 N1596 N1597 10
D1597 N1597 0 diode
R1598 N1597 N1598 10
D1598 N1598 0 diode
R1599 N1598 N1599 10
D1599 N1599 0 diode
R1600 N1599 N1600 10
D1600 N1600 0 diode
R1601 N1600 N1601 10
D1601 N1601 0 diode
R1602 N1601 N1602 10
D1602 N1602 0 diode
R1603 N1602 N1603 10
D1603 N1603 0 diode
R1604 N1603 N1604 10
D1604 N1604 0 diode
R1605 N1604 N1605 10
D1605 N1605 0 diode
R1606 N1605 N1606 10
D1606 N1606 0 diode
R1607 N1606 N1607 10
D1607 N1607 0 diode
R1608 N1607 N1608 10
D1608 N1608 0 diode
R1609 N1608 N1609 10
D1609 N1609 0 diode
R1610 N1609 N1610 10
D1610 N1610 0 diode
R1611 N1610 N1611 10
D1611 N1611 0 diode
R1612 N1611 N1612 10
D1612 N1612 0 diode
R1613 N1612 N1613 10
D1613 N1613 0 diode
R1614 N1613 N1614 10
D1614 N1614 0 diode
R1615 N1614 N1615 10
D1615 N1615 0 diode
R1616 N1615 N1616 10
D1616 N1616 0 diode
R1617 N1616 N1617 10
D1617 N1617 0 diode
R1618 N1617 N1618 10
D1618 N1618 0 diode
R1619 N1618 N1619 10
D1619 N1619 0 diode
R1620 N1619 N1620 10
D1620 N1620 0 diode
R1621 N1620 N1621 10
D1621 N1621 0 diode
R1622 N1621 N1622 10
D1622 N1622 0 diode
R1623 N1622 N1623 10
D1623 N1623 0 diode
R1624 N1623 N1624 10
D1624 N1624 0 diode
R1625 N1624 N1625 10
D1625 N1625 0 diode
R1626 N1625 N1626 10
D1626 N1626 0 diode
R1627 N1626 N1627 10
D1627 N1627 0 diode
R1628 N1627 N1628 10
D1628 N1628 0 diode
R1629 N1628 N1629 10
D1629 N1629 0 diode
R1630 N1629 N1630 10
D1630 N1630 0 diode
R1631 N1630 N1631 10
D1631 N1631 0 diode
R1632 N1631 N1632 10
D1632 N1632 0 diode
R1633 N1632 N1633 10
D1633 N1633 0 diode
R1634 N1633 N1634 10
D1634 N1634 0 diode
R1635 N1634 N1635 10
D1635 N1635 0 diode
R1636 N1635 N1636 10
D1636 N1636 0 diode
R1637 N1636 N1637 10
D1637 N1637 0 diode
R1638 N1637 N1638 10
D1638 N1638 0 diode
R1639 N1638 N1639 10
D1639 N1639 0 diode
R1640 N1639 N1640 10
D1640 N1640 0 diode
R1641 N1640 N1641 10
D1641 N1641 0 diode
R1642 N1641 N1642 10
D1642 N1642 0 diode
R1643 N1642 N1643 10
D1643 N1643 0 diode
R1644 N1643 N1644 10
D1644 N1644 0 diode
R1645 N1644 N1645 10
D1645 N1645 0 diode
R1646 N1645 N1646 10
D1646 N1646 0 diode
R1647 N1646 N1647 10
D1647 N1647 0 diode
R1648 N1647 N1648 10
D1648 N1648 0 diode
R1649 N1648 N1649 10
D1649 N1649 0 diode
R1650 N1649 N1650 10
D1650 N1650 0 diode
R1651 N1650 N1651 10
D1651 N1651 0 diode
R1652 N1651 N1652 10
D1652 N1652 0 diode
R1653 N1652 N1653 10
D1653 N1653 0 diode
R1654 N1653 N1654 10
D1654 N1654 0 diode
R1655 N1654 N1655 10
D1655 N1655 0 diode
R1656 N1655 N1656 10
D1656 N1656 0 diode
R1657 N1656 N1657 10
D1657 N1657 0 diode
R1658 N1657 N1658 10
D1658 N1658 0 diode
R1659 N1658 N1659 10
D1659 N1659 0 diode
R1660 N1659 N1660 10
D1660 N1660 0 diode
R1661 N1660 N1661 10
D1661 N1661 0 diode
R1662 N1661 N1662 10
D1662 N1662 0 diode
R1663 N1662 N1663 10
D1663 N1663 0 diode
R1664 N1663 N1664 10
D1664 N1664 0 diode
R1665 N1664 N1665 10
D1665 N1665 0 diode
R1666 N1665 N1666 10
D1666 N1666 0 diode
R1667 N1666 N1667 10
D1667 N1667 0 diode
R1668 N1667 N1668 10
D1668 N1668 0 diode
R1669 N1668 N1669 10
D1669 N1669 0 diode
R1670 N1669 N1670 10
D1670 N1670 0 diode
R1671 N1670 N1671 10
D1671 N1671 0 diode
R1672 N1671 N1672 10
D1672 N1672 0 diode
R1673 N1672 N1673 10
D1673 N1673 0 diode
R1674 N1673 N1674 10
D1674 N1674 0 diode
R1675 N1674 N1675 10
D1675 N1675 0 diode
R1676 N1675 N1676 10
D1676 N1676 0 diode
R1677 N1676 N1677 10
D1677 N1677 0 diode
R1678 N1677 N1678 10
D1678 N1678 0 diode
R1679 N1678 N1679 10
D1679 N1679 0 diode
R1680 N1679 N1680 10
D1680 N1680 0 diode
R1681 N1680 N1681 10
D1681 N1681 0 diode
R1682 N1681 N1682 10
D1682 N1682 0 diode
R1683 N1682 N1683 10
D1683 N1683 0 diode
R1684 N1683 N1684 10
D1684 N1684 0 diode
R1685 N1684 N1685 10
D1685 N1685 0 diode
R1686 N1685 N1686 10
D1686 N1686 0 diode
R1687 N1686 N1687 10
D1687 N1687 0 diode
R1688 N1687 N1688 10
D1688 N1688 0 diode
R1689 N1688 N1689 10
D1689 N1689 0 diode
R1690 N1689 N1690 10
D1690 N1690 0 diode
R1691 N1690 N1691 10
D1691 N1691 0 diode
R1692 N1691 N1692 10
D1692 N1692 0 diode
R1693 N1692 N1693 10
D1693 N1693 0 diode
R1694 N1693 N1694 10
D1694 N1694 0 diode
R1695 N1694 N1695 10
D1695 N1695 0 diode
R1696 N1695 N1696 10
D1696 N1696 0 diode
R1697 N1696 N1697 10
D1697 N1697 0 diode
R1698 N1697 N1698 10
D1698 N1698 0 diode
R1699 N1698 N1699 10
D1699 N1699 0 diode
R1700 N1699 N1700 10
D1700 N1700 0 diode
R1701 N1700 N1701 10
D1701 N1701 0 diode
R1702 N1701 N1702 10
D1702 N1702 0 diode
R1703 N1702 N1703 10
D1703 N1703 0 diode
R1704 N1703 N1704 10
D1704 N1704 0 diode
R1705 N1704 N1705 10
D1705 N1705 0 diode
R1706 N1705 N1706 10
D1706 N1706 0 diode
R1707 N1706 N1707 10
D1707 N1707 0 diode
R1708 N1707 N1708 10
D1708 N1708 0 diode
R1709 N1708 N1709 10
D1709 N1709 0 diode
R1710 N1709 N1710 10
D1710 N1710 0 diode
R1711 N1710 N1711 10
D1711 N1711 0 diode
R1712 N1711 N1712 10
D1712 N1712 0 diode
R1713 N1712 N1713 10
D1713 N1713 0 diode
R1714 N1713 N1714 10
D1714 N1714 0 diode
R1715 N1714 N1715 10
D1715 N1715 0 diode
R1716 N1715 N1716 10
D1716 N1716 0 diode
R1717 N1716 N1717 10
D1717 N1717 0 diode
R1718 N1717 N1718 10
D1718 N1718 0 diode
R1719 N1718 N1719 10
D1719 N1719 0 diode
R1720 N1719 N1720 10
D1720 N1720 0 diode
R1721 N1720 N1721 10
D1721 N1721 0 diode
R1722 N1721 N1722 10
D1722 N1722 0 diode
R1723 N1722 N1723 10
D1723 N1723 0 diode
R1724 N1723 N1724 10
D1724 N1724 0 diode
R1725 N1724 N1725 10
D1725 N1725 0 diode
R1726 N1725 N1726 10
D1726 N1726 0 diode
R1727 N1726 N1727 10
D1727 N1727 0 diode
R1728 N1727 N1728 10
D1728 N1728 0 diode
R1729 N1728 N1729 10
D1729 N1729 0 diode
R1730 N1729 N1730 10
D1730 N1730 0 diode
R1731 N1730 N1731 10
D1731 N1731 0 diode
R1732 N1731 N1732 10
D1732 N1732 0 diode
R1733 N1732 N1733 10
D1733 N1733 0 diode
R1734 N1733 N1734 10
D1734 N1734 0 diode
R1735 N1734 N1735 10
D1735 N1735 0 diode
R1736 N1735 N1736 10
D1736 N1736 0 diode
R1737 N1736 N1737 10
D1737 N1737 0 diode
R1738 N1737 N1738 10
D1738 N1738 0 diode
R1739 N1738 N1739 10
D1739 N1739 0 diode
R1740 N1739 N1740 10
D1740 N1740 0 diode
R1741 N1740 N1741 10
D1741 N1741 0 diode
R1742 N1741 N1742 10
D1742 N1742 0 diode
R1743 N1742 N1743 10
D1743 N1743 0 diode
R1744 N1743 N1744 10
D1744 N1744 0 diode
R1745 N1744 N1745 10
D1745 N1745 0 diode
R1746 N1745 N1746 10
D1746 N1746 0 diode
R1747 N1746 N1747 10
D1747 N1747 0 diode
R1748 N1747 N1748 10
D1748 N1748 0 diode
R1749 N1748 N1749 10
D1749 N1749 0 diode
R1750 N1749 N1750 10
D1750 N1750 0 diode
R1751 N1750 N1751 10
D1751 N1751 0 diode
R1752 N1751 N1752 10
D1752 N1752 0 diode
R1753 N1752 N1753 10
D1753 N1753 0 diode
R1754 N1753 N1754 10
D1754 N1754 0 diode
R1755 N1754 N1755 10
D1755 N1755 0 diode
R1756 N1755 N1756 10
D1756 N1756 0 diode
R1757 N1756 N1757 10
D1757 N1757 0 diode
R1758 N1757 N1758 10
D1758 N1758 0 diode
R1759 N1758 N1759 10
D1759 N1759 0 diode
R1760 N1759 N1760 10
D1760 N1760 0 diode
R1761 N1760 N1761 10
D1761 N1761 0 diode
R1762 N1761 N1762 10
D1762 N1762 0 diode
R1763 N1762 N1763 10
D1763 N1763 0 diode
R1764 N1763 N1764 10
D1764 N1764 0 diode
R1765 N1764 N1765 10
D1765 N1765 0 diode
R1766 N1765 N1766 10
D1766 N1766 0 diode
R1767 N1766 N1767 10
D1767 N1767 0 diode
R1768 N1767 N1768 10
D1768 N1768 0 diode
R1769 N1768 N1769 10
D1769 N1769 0 diode
R1770 N1769 N1770 10
D1770 N1770 0 diode
R1771 N1770 N1771 10
D1771 N1771 0 diode
R1772 N1771 N1772 10
D1772 N1772 0 diode
R1773 N1772 N1773 10
D1773 N1773 0 diode
R1774 N1773 N1774 10
D1774 N1774 0 diode
R1775 N1774 N1775 10
D1775 N1775 0 diode
R1776 N1775 N1776 10
D1776 N1776 0 diode
R1777 N1776 N1777 10
D1777 N1777 0 diode
R1778 N1777 N1778 10
D1778 N1778 0 diode
R1779 N1778 N1779 10
D1779 N1779 0 diode
R1780 N1779 N1780 10
D1780 N1780 0 diode
R1781 N1780 N1781 10
D1781 N1781 0 diode
R1782 N1781 N1782 10
D1782 N1782 0 diode
R1783 N1782 N1783 10
D1783 N1783 0 diode
R1784 N1783 N1784 10
D1784 N1784 0 diode
R1785 N1784 N1785 10
D1785 N1785 0 diode
R1786 N1785 N1786 10
D1786 N1786 0 diode
R1787 N1786 N1787 10
D1787 N1787 0 diode
R1788 N1787 N1788 10
D1788 N1788 0 diode
R1789 N1788 N1789 10
D1789 N1789 0 diode
R1790 N1789 N1790 10
D1790 N1790 0 diode
R1791 N1790 N1791 10
D1791 N1791 0 diode
R1792 N1791 N1792 10
D1792 N1792 0 diode
R1793 N1792 N1793 10
D1793 N1793 0 diode
R1794 N1793 N1794 10
D1794 N1794 0 diode
R1795 N1794 N1795 10
D1795 N1795 0 diode
R1796 N1795 N1796 10
D1796 N1796 0 diode
R1797 N1796 N1797 10
D1797 N1797 0 diode
R1798 N1797 N1798 10
D1798 N1798 0 diode
R1799 N1798 N1799 10
D1799 N1799 0 diode
R1800 N1799 N1800 10
D1800 N1800 0 diode
R1801 N1800 N1801 10
D1801 N1801 0 diode
R1802 N1801 N1802 10
D1802 N1802 0 diode
R1803 N1802 N1803 10
D1803 N1803 0 diode
R1804 N1803 N1804 10
D1804 N1804 0 diode
R1805 N1804 N1805 10
D1805 N1805 0 diode
R1806 N1805 N1806 10
D1806 N1806 0 diode
R1807 N1806 N1807 10
D1807 N1807 0 diode
R1808 N1807 N1808 10
D1808 N1808 0 diode
R1809 N1808 N1809 10
D1809 N1809 0 diode
R1810 N1809 N1810 10
D1810 N1810 0 diode
R1811 N1810 N1811 10
D1811 N1811 0 diode
R1812 N1811 N1812 10
D1812 N1812 0 diode
R1813 N1812 N1813 10
D1813 N1813 0 diode
R1814 N1813 N1814 10
D1814 N1814 0 diode
R1815 N1814 N1815 10
D1815 N1815 0 diode
R1816 N1815 N1816 10
D1816 N1816 0 diode
R1817 N1816 N1817 10
D1817 N1817 0 diode
R1818 N1817 N1818 10
D1818 N1818 0 diode
R1819 N1818 N1819 10
D1819 N1819 0 diode
R1820 N1819 N1820 10
D1820 N1820 0 diode
R1821 N1820 N1821 10
D1821 N1821 0 diode
R1822 N1821 N1822 10
D1822 N1822 0 diode
R1823 N1822 N1823 10
D1823 N1823 0 diode
R1824 N1823 N1824 10
D1824 N1824 0 diode
R1825 N1824 N1825 10
D1825 N1825 0 diode
R1826 N1825 N1826 10
D1826 N1826 0 diode
R1827 N1826 N1827 10
D1827 N1827 0 diode
R1828 N1827 N1828 10
D1828 N1828 0 diode
R1829 N1828 N1829 10
D1829 N1829 0 diode
R1830 N1829 N1830 10
D1830 N1830 0 diode
R1831 N1830 N1831 10
D1831 N1831 0 diode
R1832 N1831 N1832 10
D1832 N1832 0 diode
R1833 N1832 N1833 10
D1833 N1833 0 diode
R1834 N1833 N1834 10
D1834 N1834 0 diode
R1835 N1834 N1835 10
D1835 N1835 0 diode
R1836 N1835 N1836 10
D1836 N1836 0 diode
R1837 N1836 N1837 10
D1837 N1837 0 diode
R1838 N1837 N1838 10
D1838 N1838 0 diode
R1839 N1838 N1839 10
D1839 N1839 0 diode
R1840 N1839 N1840 10
D1840 N1840 0 diode
R1841 N1840 N1841 10
D1841 N1841 0 diode
R1842 N1841 N1842 10
D1842 N1842 0 diode
R1843 N1842 N1843 10
D1843 N1843 0 diode
R1844 N1843 N1844 10
D1844 N1844 0 diode
R1845 N1844 N1845 10
D1845 N1845 0 diode
R1846 N1845 N1846 10
D1846 N1846 0 diode
R1847 N1846 N1847 10
D1847 N1847 0 diode
R1848 N1847 N1848 10
D1848 N1848 0 diode
R1849 N1848 N1849 10
D1849 N1849 0 diode
R1850 N1849 N1850 10
D1850 N1850 0 diode
R1851 N1850 N1851 10
D1851 N1851 0 diode
R1852 N1851 N1852 10
D1852 N1852 0 diode
R1853 N1852 N1853 10
D1853 N1853 0 diode
R1854 N1853 N1854 10
D1854 N1854 0 diode
R1855 N1854 N1855 10
D1855 N1855 0 diode
R1856 N1855 N1856 10
D1856 N1856 0 diode
R1857 N1856 N1857 10
D1857 N1857 0 diode
R1858 N1857 N1858 10
D1858 N1858 0 diode
R1859 N1858 N1859 10
D1859 N1859 0 diode
R1860 N1859 N1860 10
D1860 N1860 0 diode
R1861 N1860 N1861 10
D1861 N1861 0 diode
R1862 N1861 N1862 10
D1862 N1862 0 diode
R1863 N1862 N1863 10
D1863 N1863 0 diode
R1864 N1863 N1864 10
D1864 N1864 0 diode
R1865 N1864 N1865 10
D1865 N1865 0 diode
R1866 N1865 N1866 10
D1866 N1866 0 diode
R1867 N1866 N1867 10
D1867 N1867 0 diode
R1868 N1867 N1868 10
D1868 N1868 0 diode
R1869 N1868 N1869 10
D1869 N1869 0 diode
R1870 N1869 N1870 10
D1870 N1870 0 diode
R1871 N1870 N1871 10
D1871 N1871 0 diode
R1872 N1871 N1872 10
D1872 N1872 0 diode
R1873 N1872 N1873 10
D1873 N1873 0 diode
R1874 N1873 N1874 10
D1874 N1874 0 diode
R1875 N1874 N1875 10
D1875 N1875 0 diode
R1876 N1875 N1876 10
D1876 N1876 0 diode
R1877 N1876 N1877 10
D1877 N1877 0 diode
R1878 N1877 N1878 10
D1878 N1878 0 diode
R1879 N1878 N1879 10
D1879 N1879 0 diode
R1880 N1879 N1880 10
D1880 N1880 0 diode
R1881 N1880 N1881 10
D1881 N1881 0 diode
R1882 N1881 N1882 10
D1882 N1882 0 diode
R1883 N1882 N1883 10
D1883 N1883 0 diode
R1884 N1883 N1884 10
D1884 N1884 0 diode
R1885 N1884 N1885 10
D1885 N1885 0 diode
R1886 N1885 N1886 10
D1886 N1886 0 diode
R1887 N1886 N1887 10
D1887 N1887 0 diode
R1888 N1887 N1888 10
D1888 N1888 0 diode
R1889 N1888 N1889 10
D1889 N1889 0 diode
R1890 N1889 N1890 10
D1890 N1890 0 diode
R1891 N1890 N1891 10
D1891 N1891 0 diode
R1892 N1891 N1892 10
D1892 N1892 0 diode
R1893 N1892 N1893 10
D1893 N1893 0 diode
R1894 N1893 N1894 10
D1894 N1894 0 diode
R1895 N1894 N1895 10
D1895 N1895 0 diode
R1896 N1895 N1896 10
D1896 N1896 0 diode
R1897 N1896 N1897 10
D1897 N1897 0 diode
R1898 N1897 N1898 10
D1898 N1898 0 diode
R1899 N1898 N1899 10
D1899 N1899 0 diode
R1900 N1899 N1900 10
D1900 N1900 0 diode
R1901 N1900 N1901 10
D1901 N1901 0 diode
R1902 N1901 N1902 10
D1902 N1902 0 diode
R1903 N1902 N1903 10
D1903 N1903 0 diode
R1904 N1903 N1904 10
D1904 N1904 0 diode
R1905 N1904 N1905 10
D1905 N1905 0 diode
R1906 N1905 N1906 10
D1906 N1906 0 diode
R1907 N1906 N1907 10
D1907 N1907 0 diode
R1908 N1907 N1908 10
D1908 N1908 0 diode
R1909 N1908 N1909 10
D1909 N1909 0 diode
R1910 N1909 N1910 10
D1910 N1910 0 diode
R1911 N1910 N1911 10
D1911 N1911 0 diode
R1912 N1911 N1912 10
D1912 N1912 0 diode
R1913 N1912 N1913 10
D1913 N1913 0 diode
R1914 N1913 N1914 10
D1914 N1914 0 diode
R1915 N1914 N1915 10
D1915 N1915 0 diode
R1916 N1915 N1916 10
D1916 N1916 0 diode
R1917 N1916 N1917 10
D1917 N1917 0 diode
R1918 N1917 N1918 10
D1918 N1918 0 diode
R1919 N1918 N1919 10
D1919 N1919 0 diode
R1920 N1919 N1920 10
D1920 N1920 0 diode
R1921 N1920 N1921 10
D1921 N1921 0 diode
R1922 N1921 N1922 10
D1922 N1922 0 diode
R1923 N1922 N1923 10
D1923 N1923 0 diode
R1924 N1923 N1924 10
D1924 N1924 0 diode
R1925 N1924 N1925 10
D1925 N1925 0 diode
R1926 N1925 N1926 10
D1926 N1926 0 diode
R1927 N1926 N1927 10
D1927 N1927 0 diode
R1928 N1927 N1928 10
D1928 N1928 0 diode
R1929 N1928 N1929 10
D1929 N1929 0 diode
R1930 N1929 N1930 10
D1930 N1930 0 diode
R1931 N1930 N1931 10
D1931 N1931 0 diode
R1932 N1931 N1932 10
D1932 N1932 0 diode
R1933 N1932 N1933 10
D1933 N1933 0 diode
R1934 N1933 N1934 10
D1934 N1934 0 diode
R1935 N1934 N1935 10
D1935 N1935 0 diode
R1936 N1935 N1936 10
D1936 N1936 0 diode
R1937 N1936 N1937 10
D1937 N1937 0 diode
R1938 N1937 N1938 10
D1938 N1938 0 diode
R1939 N1938 N1939 10
D1939 N1939 0 diode
R1940 N1939 N1940 10
D1940 N1940 0 diode
R1941 N1940 N1941 10
D1941 N1941 0 diode
R1942 N1941 N1942 10
D1942 N1942 0 diode
R1943 N1942 N1943 10
D1943 N1943 0 diode
R1944 N1943 N1944 10
D1944 N1944 0 diode
R1945 N1944 N1945 10
D1945 N1945 0 diode
R1946 N1945 N1946 10
D1946 N1946 0 diode
R1947 N1946 N1947 10
D1947 N1947 0 diode
R1948 N1947 N1948 10
D1948 N1948 0 diode
R1949 N1948 N1949 10
D1949 N1949 0 diode
R1950 N1949 N1950 10
D1950 N1950 0 diode
R1951 N1950 N1951 10
D1951 N1951 0 diode
R1952 N1951 N1952 10
D1952 N1952 0 diode
R1953 N1952 N1953 10
D1953 N1953 0 diode
R1954 N1953 N1954 10
D1954 N1954 0 diode
R1955 N1954 N1955 10
D1955 N1955 0 diode
R1956 N1955 N1956 10
D1956 N1956 0 diode
R1957 N1956 N1957 10
D1957 N1957 0 diode
R1958 N1957 N1958 10
D1958 N1958 0 diode
R1959 N1958 N1959 10
D1959 N1959 0 diode
R1960 N1959 N1960 10
D1960 N1960 0 diode
R1961 N1960 N1961 10
D1961 N1961 0 diode
R1962 N1961 N1962 10
D1962 N1962 0 diode
R1963 N1962 N1963 10
D1963 N1963 0 diode
R1964 N1963 N1964 10
D1964 N1964 0 diode
R1965 N1964 N1965 10
D1965 N1965 0 diode
R1966 N1965 N1966 10
D1966 N1966 0 diode
R1967 N1966 N1967 10
D1967 N1967 0 diode
R1968 N1967 N1968 10
D1968 N1968 0 diode
R1969 N1968 N1969 10
D1969 N1969 0 diode
R1970 N1969 N1970 10
D1970 N1970 0 diode
R1971 N1970 N1971 10
D1971 N1971 0 diode
R1972 N1971 N1972 10
D1972 N1972 0 diode
R1973 N1972 N1973 10
D1973 N1973 0 diode
R1974 N1973 N1974 10
D1974 N1974 0 diode
R1975 N1974 N1975 10
D1975 N1975 0 diode
R1976 N1975 N1976 10
D1976 N1976 0 diode
R1977 N1976 N1977 10
D1977 N1977 0 diode
R1978 N1977 N1978 10
D1978 N1978 0 diode
R1979 N1978 N1979 10
D1979 N1979 0 diode
R1980 N1979 N1980 10
D1980 N1980 0 diode
R1981 N1980 N1981 10
D1981 N1981 0 diode
R1982 N1981 N1982 10
D1982 N1982 0 diode
R1983 N1982 N1983 10
D1983 N1983 0 diode
R1984 N1983 N1984 10
D1984 N1984 0 diode
R1985 N1984 N1985 10
D1985 N1985 0 diode
R1986 N1985 N1986 10
D1986 N1986 0 diode
R1987 N1986 N1987 10
D1987 N1987 0 diode
R1988 N1987 N1988 10
D1988 N1988 0 diode
R1989 N1988 N1989 10
D1989 N1989 0 diode
R1990 N1989 N1990 10
D1990 N1990 0 diode
R1991 N1990 N1991 10
D1991 N1991 0 diode
R1992 N1991 N1992 10
D1992 N1992 0 diode
R1993 N1992 N1993 10
D1993 N1993 0 diode
R1994 N1993 N1994 10
D1994 N1994 0 diode
R1995 N1994 N1995 10
D1995 N1995 0 diode
R1996 N1995 N1996 10
D1996 N1996 0 diode
R1997 N1996 N1997 10
D1997 N1997 0 diode
R1998 N1997 N1998 10
D1998 N1998 0 diode
R1999 N1998 N1999 10
D1999 N1999 0 diode
R2000 N1999 N2000 10
D2000 N2000 0 diode
R2001 N2000 N2001 10
D2001 N2001 0 diode
R2002 N2001 N2002 10
D2002 N2002 0 diode
R2003 N2002 N2003 10
D2003 N2003 0 diode
R2004 N2003 N2004 10
D2004 N2004 0 diode
R2005 N2004 N2005 10
D2005 N2005 0 diode
R2006 N2005 N2006 10
D2006 N2006 0 diode
R2007 N2006 N2007 10
D2007 N2007 0 diode
R2008 N2007 N2008 10
D2008 N2008 0 diode
R2009 N2008 N2009 10
D2009 N2009 0 diode
R2010 N2009 N2010 10
D2010 N2010 0 diode
R2011 N2010 N2011 10
D2011 N2011 0 diode
R2012 N2011 N2012 10
D2012 N2012 0 diode
R2013 N2012 N2013 10
D2013 N2013 0 diode
R2014 N2013 N2014 10
D2014 N2014 0 diode
R2015 N2014 N2015 10
D2015 N2015 0 diode
R2016 N2015 N2016 10
D2016 N2016 0 diode
R2017 N2016 N2017 10
D2017 N2017 0 diode
R2018 N2017 N2018 10
D2018 N2018 0 diode
R2019 N2018 N2019 10
D2019 N2019 0 diode
R2020 N2019 N2020 10
D2020 N2020 0 diode
R2021 N2020 N2021 10
D2021 N2021 0 diode
R2022 N2021 N2022 10
D2022 N2022 0 diode
R2023 N2022 N2023 10
D2023 N2023 0 diode
R2024 N2023 N2024 10
D2024 N2024 0 diode
R2025 N2024 N2025 10
D2025 N2025 0 diode
R2026 N2025 N2026 10
D2026 N2026 0 diode
R2027 N2026 N2027 10
D2027 N2027 0 diode
R2028 N2027 N2028 10
D2028 N2028 0 diode
R2029 N2028 N2029 10
D2029 N2029 0 diode
R2030 N2029 N2030 10
D2030 N2030 0 diode
R2031 N2030 N2031 10
D2031 N2031 0 diode
R2032 N2031 N2032 10
D2032 N2032 0 diode
R2033 N2032 N2033 10
D2033 N2033 0 diode
R2034 N2033 N2034 10
D2034 N2034 0 diode
R2035 N2034 N2035 10
D2035 N2035 0 diode
R2036 N2035 N2036 10
D2036 N2036 0 diode
R2037 N2036 N2037 10
D2037 N2037 0 diode
R2038 N2037 N2038 10
D2038 N2038 0 diode
R2039 N2038 N2039 10
D2039 N2039 0 diode
R2040 N2039 N2040 10
D2040 N2040 0 diode
R2041 N2040 N2041 10
D2041 N2041 0 diode
R2042 N2041 N2042 10
D2042 N2042 0 diode
R2043 N2042 N2043 10
D2043 N2043 0 diode
R2044 N2043 N2044 10
D2044 N2044 0 diode
R2045 N2044 N2045 10
D2045 N2045 0 diode
R2046 N2045 N2046 10
D2046 N2046 0 diode
R2047 N2046 N2047 10
D2047 N2047 0 diode
R2048 N2047 N2048 10
D2048 N2048 0 diode
R2049 N2048 N2049 10
D2049 N2049 0 diode
R2050 N2049 N2050 10
D2050 N2050 0 diode
R2051 N2050 N2051 10
D2051 N2051 0 diode
R2052 N2051 N2052 10
D2052 N2052 0 diode
R2053 N2052 N2053 10
D2053 N2053 0 diode
R2054 N2053 N2054 10
D2054 N2054 0 diode
R2055 N2054 N2055 10
D2055 N2055 0 diode
R2056 N2055 N2056 10
D2056 N2056 0 diode
R2057 N2056 N2057 10
D2057 N2057 0 diode
R2058 N2057 N2058 10
D2058 N2058 0 diode
R2059 N2058 N2059 10
D2059 N2059 0 diode
R2060 N2059 N2060 10
D2060 N2060 0 diode
R2061 N2060 N2061 10
D2061 N2061 0 diode
R2062 N2061 N2062 10
D2062 N2062 0 diode
R2063 N2062 N2063 10
D2063 N2063 0 diode
R2064 N2063 N2064 10
D2064 N2064 0 diode
R2065 N2064 N2065 10
D2065 N2065 0 diode
R2066 N2065 N2066 10
D2066 N2066 0 diode
R2067 N2066 N2067 10
D2067 N2067 0 diode
R2068 N2067 N2068 10
D2068 N2068 0 diode
R2069 N2068 N2069 10
D2069 N2069 0 diode
R2070 N2069 N2070 10
D2070 N2070 0 diode
R2071 N2070 N2071 10
D2071 N2071 0 diode
R2072 N2071 N2072 10
D2072 N2072 0 diode
R2073 N2072 N2073 10
D2073 N2073 0 diode
R2074 N2073 N2074 10
D2074 N2074 0 diode
R2075 N2074 N2075 10
D2075 N2075 0 diode
R2076 N2075 N2076 10
D2076 N2076 0 diode
R2077 N2076 N2077 10
D2077 N2077 0 diode
R2078 N2077 N2078 10
D2078 N2078 0 diode
R2079 N2078 N2079 10
D2079 N2079 0 diode
R2080 N2079 N2080 10
D2080 N2080 0 diode
R2081 N2080 N2081 10
D2081 N2081 0 diode
R2082 N2081 N2082 10
D2082 N2082 0 diode
R2083 N2082 N2083 10
D2083 N2083 0 diode
R2084 N2083 N2084 10
D2084 N2084 0 diode
R2085 N2084 N2085 10
D2085 N2085 0 diode
R2086 N2085 N2086 10
D2086 N2086 0 diode
R2087 N2086 N2087 10
D2087 N2087 0 diode
R2088 N2087 N2088 10
D2088 N2088 0 diode
R2089 N2088 N2089 10
D2089 N2089 0 diode
R2090 N2089 N2090 10
D2090 N2090 0 diode
R2091 N2090 N2091 10
D2091 N2091 0 diode
R2092 N2091 N2092 10
D2092 N2092 0 diode
R2093 N2092 N2093 10
D2093 N2093 0 diode
R2094 N2093 N2094 10
D2094 N2094 0 diode
R2095 N2094 N2095 10
D2095 N2095 0 diode
R2096 N2095 N2096 10
D2096 N2096 0 diode
R2097 N2096 N2097 10
D2097 N2097 0 diode
R2098 N2097 N2098 10
D2098 N2098 0 diode
R2099 N2098 N2099 10
D2099 N2099 0 diode
R2100 N2099 N2100 10
D2100 N2100 0 diode
R2101 N2100 N2101 10
D2101 N2101 0 diode
R2102 N2101 N2102 10
D2102 N2102 0 diode
R2103 N2102 N2103 10
D2103 N2103 0 diode
R2104 N2103 N2104 10
D2104 N2104 0 diode
R2105 N2104 N2105 10
D2105 N2105 0 diode
R2106 N2105 N2106 10
D2106 N2106 0 diode
R2107 N2106 N2107 10
D2107 N2107 0 diode
R2108 N2107 N2108 10
D2108 N2108 0 diode
R2109 N2108 N2109 10
D2109 N2109 0 diode
R2110 N2109 N2110 10
D2110 N2110 0 diode
R2111 N2110 N2111 10
D2111 N2111 0 diode
R2112 N2111 N2112 10
D2112 N2112 0 diode
R2113 N2112 N2113 10
D2113 N2113 0 diode
R2114 N2113 N2114 10
D2114 N2114 0 diode
R2115 N2114 N2115 10
D2115 N2115 0 diode
R2116 N2115 N2116 10
D2116 N2116 0 diode
R2117 N2116 N2117 10
D2117 N2117 0 diode
R2118 N2117 N2118 10
D2118 N2118 0 diode
R2119 N2118 N2119 10
D2119 N2119 0 diode
R2120 N2119 N2120 10
D2120 N2120 0 diode
R2121 N2120 N2121 10
D2121 N2121 0 diode
R2122 N2121 N2122 10
D2122 N2122 0 diode
R2123 N2122 N2123 10
D2123 N2123 0 diode
R2124 N2123 N2124 10
D2124 N2124 0 diode
R2125 N2124 N2125 10
D2125 N2125 0 diode
R2126 N2125 N2126 10
D2126 N2126 0 diode
R2127 N2126 N2127 10
D2127 N2127 0 diode
R2128 N2127 N2128 10
D2128 N2128 0 diode
R2129 N2128 N2129 10
D2129 N2129 0 diode
R2130 N2129 N2130 10
D2130 N2130 0 diode
R2131 N2130 N2131 10
D2131 N2131 0 diode
R2132 N2131 N2132 10
D2132 N2132 0 diode
R2133 N2132 N2133 10
D2133 N2133 0 diode
R2134 N2133 N2134 10
D2134 N2134 0 diode
R2135 N2134 N2135 10
D2135 N2135 0 diode
R2136 N2135 N2136 10
D2136 N2136 0 diode
R2137 N2136 N2137 10
D2137 N2137 0 diode
R2138 N2137 N2138 10
D2138 N2138 0 diode
R2139 N2138 N2139 10
D2139 N2139 0 diode
R2140 N2139 N2140 10
D2140 N2140 0 diode
R2141 N2140 N2141 10
D2141 N2141 0 diode
R2142 N2141 N2142 10
D2142 N2142 0 diode
R2143 N2142 N2143 10
D2143 N2143 0 diode
R2144 N2143 N2144 10
D2144 N2144 0 diode
R2145 N2144 N2145 10
D2145 N2145 0 diode
R2146 N2145 N2146 10
D2146 N2146 0 diode
R2147 N2146 N2147 10
D2147 N2147 0 diode
R2148 N2147 N2148 10
D2148 N2148 0 diode
R2149 N2148 N2149 10
D2149 N2149 0 diode
R2150 N2149 N2150 10
D2150 N2150 0 diode
R2151 N2150 N2151 10
D2151 N2151 0 diode
R2152 N2151 N2152 10
D2152 N2152 0 diode
R2153 N2152 N2153 10
D2153 N2153 0 diode
R2154 N2153 N2154 10
D2154 N2154 0 diode
R2155 N2154 N2155 10
D2155 N2155 0 diode
R2156 N2155 N2156 10
D2156 N2156 0 diode
R2157 N2156 N2157 10
D2157 N2157 0 diode
R2158 N2157 N2158 10
D2158 N2158 0 diode
R2159 N2158 N2159 10
D2159 N2159 0 diode
R2160 N2159 N2160 10
D2160 N2160 0 diode
R2161 N2160 N2161 10
D2161 N2161 0 diode
R2162 N2161 N2162 10
D2162 N2162 0 diode
R2163 N2162 N2163 10
D2163 N2163 0 diode
R2164 N2163 N2164 10
D2164 N2164 0 diode
R2165 N2164 N2165 10
D2165 N2165 0 diode
R2166 N2165 N2166 10
D2166 N2166 0 diode
R2167 N2166 N2167 10
D2167 N2167 0 diode
R2168 N2167 N2168 10
D2168 N2168 0 diode
R2169 N2168 N2169 10
D2169 N2169 0 diode
R2170 N2169 N2170 10
D2170 N2170 0 diode
R2171 N2170 N2171 10
D2171 N2171 0 diode
R2172 N2171 N2172 10
D2172 N2172 0 diode
R2173 N2172 N2173 10
D2173 N2173 0 diode
R2174 N2173 N2174 10
D2174 N2174 0 diode
R2175 N2174 N2175 10
D2175 N2175 0 diode
R2176 N2175 N2176 10
D2176 N2176 0 diode
R2177 N2176 N2177 10
D2177 N2177 0 diode
R2178 N2177 N2178 10
D2178 N2178 0 diode
R2179 N2178 N2179 10
D2179 N2179 0 diode
R2180 N2179 N2180 10
D2180 N2180 0 diode
R2181 N2180 N2181 10
D2181 N2181 0 diode
R2182 N2181 N2182 10
D2182 N2182 0 diode
R2183 N2182 N2183 10
D2183 N2183 0 diode
R2184 N2183 N2184 10
D2184 N2184 0 diode
R2185 N2184 N2185 10
D2185 N2185 0 diode
R2186 N2185 N2186 10
D2186 N2186 0 diode
R2187 N2186 N2187 10
D2187 N2187 0 diode
R2188 N2187 N2188 10
D2188 N2188 0 diode
R2189 N2188 N2189 10
D2189 N2189 0 diode
R2190 N2189 N2190 10
D2190 N2190 0 diode
R2191 N2190 N2191 10
D2191 N2191 0 diode
R2192 N2191 N2192 10
D2192 N2192 0 diode
R2193 N2192 N2193 10
D2193 N2193 0 diode
R2194 N2193 N2194 10
D2194 N2194 0 diode
R2195 N2194 N2195 10
D2195 N2195 0 diode
R2196 N2195 N2196 10
D2196 N2196 0 diode
R2197 N2196 N2197 10
D2197 N2197 0 diode
R2198 N2197 N2198 10
D2198 N2198 0 diode
R2199 N2198 N2199 10
D2199 N2199 0 diode
R2200 N2199 N2200 10
D2200 N2200 0 diode
R2201 N2200 N2201 10
D2201 N2201 0 diode
R2202 N2201 N2202 10
D2202 N2202 0 diode
R2203 N2202 N2203 10
D2203 N2203 0 diode
R2204 N2203 N2204 10
D2204 N2204 0 diode
R2205 N2204 N2205 10
D2205 N2205 0 diode
R2206 N2205 N2206 10
D2206 N2206 0 diode
R2207 N2206 N2207 10
D2207 N2207 0 diode
R2208 N2207 N2208 10
D2208 N2208 0 diode
R2209 N2208 N2209 10
D2209 N2209 0 diode
R2210 N2209 N2210 10
D2210 N2210 0 diode
R2211 N2210 N2211 10
D2211 N2211 0 diode
R2212 N2211 N2212 10
D2212 N2212 0 diode
R2213 N2212 N2213 10
D2213 N2213 0 diode
R2214 N2213 N2214 10
D2214 N2214 0 diode
R2215 N2214 N2215 10
D2215 N2215 0 diode
R2216 N2215 N2216 10
D2216 N2216 0 diode
R2217 N2216 N2217 10
D2217 N2217 0 diode
R2218 N2217 N2218 10
D2218 N2218 0 diode
R2219 N2218 N2219 10
D2219 N2219 0 diode
R2220 N2219 N2220 10
D2220 N2220 0 diode
R2221 N2220 N2221 10
D2221 N2221 0 diode
R2222 N2221 N2222 10
D2222 N2222 0 diode
R2223 N2222 N2223 10
D2223 N2223 0 diode
R2224 N2223 N2224 10
D2224 N2224 0 diode
R2225 N2224 N2225 10
D2225 N2225 0 diode
R2226 N2225 N2226 10
D2226 N2226 0 diode
R2227 N2226 N2227 10
D2227 N2227 0 diode
R2228 N2227 N2228 10
D2228 N2228 0 diode
R2229 N2228 N2229 10
D2229 N2229 0 diode
R2230 N2229 N2230 10
D2230 N2230 0 diode
R2231 N2230 N2231 10
D2231 N2231 0 diode
R2232 N2231 N2232 10
D2232 N2232 0 diode
R2233 N2232 N2233 10
D2233 N2233 0 diode
R2234 N2233 N2234 10
D2234 N2234 0 diode
R2235 N2234 N2235 10
D2235 N2235 0 diode
R2236 N2235 N2236 10
D2236 N2236 0 diode
R2237 N2236 N2237 10
D2237 N2237 0 diode
R2238 N2237 N2238 10
D2238 N2238 0 diode
R2239 N2238 N2239 10
D2239 N2239 0 diode
R2240 N2239 N2240 10
D2240 N2240 0 diode
R2241 N2240 N2241 10
D2241 N2241 0 diode
R2242 N2241 N2242 10
D2242 N2242 0 diode
R2243 N2242 N2243 10
D2243 N2243 0 diode
R2244 N2243 N2244 10
D2244 N2244 0 diode
R2245 N2244 N2245 10
D2245 N2245 0 diode
R2246 N2245 N2246 10
D2246 N2246 0 diode
R2247 N2246 N2247 10
D2247 N2247 0 diode
R2248 N2247 N2248 10
D2248 N2248 0 diode
R2249 N2248 N2249 10
D2249 N2249 0 diode
R2250 N2249 N2250 10
D2250 N2250 0 diode
R2251 N2250 N2251 10
D2251 N2251 0 diode
R2252 N2251 N2252 10
D2252 N2252 0 diode
R2253 N2252 N2253 10
D2253 N2253 0 diode
R2254 N2253 N2254 10
D2254 N2254 0 diode
R2255 N2254 N2255 10
D2255 N2255 0 diode
R2256 N2255 N2256 10
D2256 N2256 0 diode
R2257 N2256 N2257 10
D2257 N2257 0 diode
R2258 N2257 N2258 10
D2258 N2258 0 diode
R2259 N2258 N2259 10
D2259 N2259 0 diode
R2260 N2259 N2260 10
D2260 N2260 0 diode
R2261 N2260 N2261 10
D2261 N2261 0 diode
R2262 N2261 N2262 10
D2262 N2262 0 diode
R2263 N2262 N2263 10
D2263 N2263 0 diode
R2264 N2263 N2264 10
D2264 N2264 0 diode
R2265 N2264 N2265 10
D2265 N2265 0 diode
R2266 N2265 N2266 10
D2266 N2266 0 diode
R2267 N2266 N2267 10
D2267 N2267 0 diode
R2268 N2267 N2268 10
D2268 N2268 0 diode
R2269 N2268 N2269 10
D2269 N2269 0 diode
R2270 N2269 N2270 10
D2270 N2270 0 diode
R2271 N2270 N2271 10
D2271 N2271 0 diode
R2272 N2271 N2272 10
D2272 N2272 0 diode
R2273 N2272 N2273 10
D2273 N2273 0 diode
R2274 N2273 N2274 10
D2274 N2274 0 diode
R2275 N2274 N2275 10
D2275 N2275 0 diode
R2276 N2275 N2276 10
D2276 N2276 0 diode
R2277 N2276 N2277 10
D2277 N2277 0 diode
R2278 N2277 N2278 10
D2278 N2278 0 diode
R2279 N2278 N2279 10
D2279 N2279 0 diode
R2280 N2279 N2280 10
D2280 N2280 0 diode
R2281 N2280 N2281 10
D2281 N2281 0 diode
R2282 N2281 N2282 10
D2282 N2282 0 diode
R2283 N2282 N2283 10
D2283 N2283 0 diode
R2284 N2283 N2284 10
D2284 N2284 0 diode
R2285 N2284 N2285 10
D2285 N2285 0 diode
R2286 N2285 N2286 10
D2286 N2286 0 diode
R2287 N2286 N2287 10
D2287 N2287 0 diode
R2288 N2287 N2288 10
D2288 N2288 0 diode
R2289 N2288 N2289 10
D2289 N2289 0 diode
R2290 N2289 N2290 10
D2290 N2290 0 diode
R2291 N2290 N2291 10
D2291 N2291 0 diode
R2292 N2291 N2292 10
D2292 N2292 0 diode
R2293 N2292 N2293 10
D2293 N2293 0 diode
R2294 N2293 N2294 10
D2294 N2294 0 diode
R2295 N2294 N2295 10
D2295 N2295 0 diode
R2296 N2295 N2296 10
D2296 N2296 0 diode
R2297 N2296 N2297 10
D2297 N2297 0 diode
R2298 N2297 N2298 10
D2298 N2298 0 diode
R2299 N2298 N2299 10
D2299 N2299 0 diode
R2300 N2299 N2300 10
D2300 N2300 0 diode
R2301 N2300 N2301 10
D2301 N2301 0 diode
R2302 N2301 N2302 10
D2302 N2302 0 diode
R2303 N2302 N2303 10
D2303 N2303 0 diode
R2304 N2303 N2304 10
D2304 N2304 0 diode
R2305 N2304 N2305 10
D2305 N2305 0 diode
R2306 N2305 N2306 10
D2306 N2306 0 diode
R2307 N2306 N2307 10
D2307 N2307 0 diode
R2308 N2307 N2308 10
D2308 N2308 0 diode
R2309 N2308 N2309 10
D2309 N2309 0 diode
R2310 N2309 N2310 10
D2310 N2310 0 diode
R2311 N2310 N2311 10
D2311 N2311 0 diode
R2312 N2311 N2312 10
D2312 N2312 0 diode
R2313 N2312 N2313 10
D2313 N2313 0 diode
R2314 N2313 N2314 10
D2314 N2314 0 diode
R2315 N2314 N2315 10
D2315 N2315 0 diode
R2316 N2315 N2316 10
D2316 N2316 0 diode
R2317 N2316 N2317 10
D2317 N2317 0 diode
R2318 N2317 N2318 10
D2318 N2318 0 diode
R2319 N2318 N2319 10
D2319 N2319 0 diode
R2320 N2319 N2320 10
D2320 N2320 0 diode
R2321 N2320 N2321 10
D2321 N2321 0 diode
R2322 N2321 N2322 10
D2322 N2322 0 diode
R2323 N2322 N2323 10
D2323 N2323 0 diode
R2324 N2323 N2324 10
D2324 N2324 0 diode
R2325 N2324 N2325 10
D2325 N2325 0 diode
R2326 N2325 N2326 10
D2326 N2326 0 diode
R2327 N2326 N2327 10
D2327 N2327 0 diode
R2328 N2327 N2328 10
D2328 N2328 0 diode
R2329 N2328 N2329 10
D2329 N2329 0 diode
R2330 N2329 N2330 10
D2330 N2330 0 diode
R2331 N2330 N2331 10
D2331 N2331 0 diode
R2332 N2331 N2332 10
D2332 N2332 0 diode
R2333 N2332 N2333 10
D2333 N2333 0 diode
R2334 N2333 N2334 10
D2334 N2334 0 diode
R2335 N2334 N2335 10
D2335 N2335 0 diode
R2336 N2335 N2336 10
D2336 N2336 0 diode
R2337 N2336 N2337 10
D2337 N2337 0 diode
R2338 N2337 N2338 10
D2338 N2338 0 diode
R2339 N2338 N2339 10
D2339 N2339 0 diode
R2340 N2339 N2340 10
D2340 N2340 0 diode
R2341 N2340 N2341 10
D2341 N2341 0 diode
R2342 N2341 N2342 10
D2342 N2342 0 diode
R2343 N2342 N2343 10
D2343 N2343 0 diode
R2344 N2343 N2344 10
D2344 N2344 0 diode
R2345 N2344 N2345 10
D2345 N2345 0 diode
R2346 N2345 N2346 10
D2346 N2346 0 diode
R2347 N2346 N2347 10
D2347 N2347 0 diode
R2348 N2347 N2348 10
D2348 N2348 0 diode
R2349 N2348 N2349 10
D2349 N2349 0 diode
R2350 N2349 N2350 10
D2350 N2350 0 diode
R2351 N2350 N2351 10
D2351 N2351 0 diode
R2352 N2351 N2352 10
D2352 N2352 0 diode
R2353 N2352 N2353 10
D2353 N2353 0 diode
R2354 N2353 N2354 10
D2354 N2354 0 diode
R2355 N2354 N2355 10
D2355 N2355 0 diode
R2356 N2355 N2356 10
D2356 N2356 0 diode
R2357 N2356 N2357 10
D2357 N2357 0 diode
R2358 N2357 N2358 10
D2358 N2358 0 diode
R2359 N2358 N2359 10
D2359 N2359 0 diode
R2360 N2359 N2360 10
D2360 N2360 0 diode
R2361 N2360 N2361 10
D2361 N2361 0 diode
R2362 N2361 N2362 10
D2362 N2362 0 diode
R2363 N2362 N2363 10
D2363 N2363 0 diode
R2364 N2363 N2364 10
D2364 N2364 0 diode
R2365 N2364 N2365 10
D2365 N2365 0 diode
R2366 N2365 N2366 10
D2366 N2366 0 diode
R2367 N2366 N2367 10
D2367 N2367 0 diode
R2368 N2367 N2368 10
D2368 N2368 0 diode
R2369 N2368 N2369 10
D2369 N2369 0 diode
R2370 N2369 N2370 10
D2370 N2370 0 diode
R2371 N2370 N2371 10
D2371 N2371 0 diode
R2372 N2371 N2372 10
D2372 N2372 0 diode
R2373 N2372 N2373 10
D2373 N2373 0 diode
R2374 N2373 N2374 10
D2374 N2374 0 diode
R2375 N2374 N2375 10
D2375 N2375 0 diode
R2376 N2375 N2376 10
D2376 N2376 0 diode
R2377 N2376 N2377 10
D2377 N2377 0 diode
R2378 N2377 N2378 10
D2378 N2378 0 diode
R2379 N2378 N2379 10
D2379 N2379 0 diode
R2380 N2379 N2380 10
D2380 N2380 0 diode
R2381 N2380 N2381 10
D2381 N2381 0 diode
R2382 N2381 N2382 10
D2382 N2382 0 diode
R2383 N2382 N2383 10
D2383 N2383 0 diode
R2384 N2383 N2384 10
D2384 N2384 0 diode
R2385 N2384 N2385 10
D2385 N2385 0 diode
R2386 N2385 N2386 10
D2386 N2386 0 diode
R2387 N2386 N2387 10
D2387 N2387 0 diode
R2388 N2387 N2388 10
D2388 N2388 0 diode
R2389 N2388 N2389 10
D2389 N2389 0 diode
R2390 N2389 N2390 10
D2390 N2390 0 diode
R2391 N2390 N2391 10
D2391 N2391 0 diode
R2392 N2391 N2392 10
D2392 N2392 0 diode
R2393 N2392 N2393 10
D2393 N2393 0 diode
R2394 N2393 N2394 10
D2394 N2394 0 diode
R2395 N2394 N2395 10
D2395 N2395 0 diode
R2396 N2395 N2396 10
D2396 N2396 0 diode
R2397 N2396 N2397 10
D2397 N2397 0 diode
R2398 N2397 N2398 10
D2398 N2398 0 diode
R2399 N2398 N2399 10
D2399 N2399 0 diode
R2400 N2399 N2400 10
D2400 N2400 0 diode
R2401 N2400 N2401 10
D2401 N2401 0 diode
R2402 N2401 N2402 10
D2402 N2402 0 diode
R2403 N2402 N2403 10
D2403 N2403 0 diode
R2404 N2403 N2404 10
D2404 N2404 0 diode
R2405 N2404 N2405 10
D2405 N2405 0 diode
R2406 N2405 N2406 10
D2406 N2406 0 diode
R2407 N2406 N2407 10
D2407 N2407 0 diode
R2408 N2407 N2408 10
D2408 N2408 0 diode
R2409 N2408 N2409 10
D2409 N2409 0 diode
R2410 N2409 N2410 10
D2410 N2410 0 diode
R2411 N2410 N2411 10
D2411 N2411 0 diode
R2412 N2411 N2412 10
D2412 N2412 0 diode
R2413 N2412 N2413 10
D2413 N2413 0 diode
R2414 N2413 N2414 10
D2414 N2414 0 diode
R2415 N2414 N2415 10
D2415 N2415 0 diode
R2416 N2415 N2416 10
D2416 N2416 0 diode
R2417 N2416 N2417 10
D2417 N2417 0 diode
R2418 N2417 N2418 10
D2418 N2418 0 diode
R2419 N2418 N2419 10
D2419 N2419 0 diode
R2420 N2419 N2420 10
D2420 N2420 0 diode
R2421 N2420 N2421 10
D2421 N2421 0 diode
R2422 N2421 N2422 10
D2422 N2422 0 diode
R2423 N2422 N2423 10
D2423 N2423 0 diode
R2424 N2423 N2424 10
D2424 N2424 0 diode
R2425 N2424 N2425 10
D2425 N2425 0 diode
R2426 N2425 N2426 10
D2426 N2426 0 diode
R2427 N2426 N2427 10
D2427 N2427 0 diode
R2428 N2427 N2428 10
D2428 N2428 0 diode
R2429 N2428 N2429 10
D2429 N2429 0 diode
R2430 N2429 N2430 10
D2430 N2430 0 diode
R2431 N2430 N2431 10
D2431 N2431 0 diode
R2432 N2431 N2432 10
D2432 N2432 0 diode
R2433 N2432 N2433 10
D2433 N2433 0 diode
R2434 N2433 N2434 10
D2434 N2434 0 diode
R2435 N2434 N2435 10
D2435 N2435 0 diode
R2436 N2435 N2436 10
D2436 N2436 0 diode
R2437 N2436 N2437 10
D2437 N2437 0 diode
R2438 N2437 N2438 10
D2438 N2438 0 diode
R2439 N2438 N2439 10
D2439 N2439 0 diode
R2440 N2439 N2440 10
D2440 N2440 0 diode
R2441 N2440 N2441 10
D2441 N2441 0 diode
R2442 N2441 N2442 10
D2442 N2442 0 diode
R2443 N2442 N2443 10
D2443 N2443 0 diode
R2444 N2443 N2444 10
D2444 N2444 0 diode
R2445 N2444 N2445 10
D2445 N2445 0 diode
R2446 N2445 N2446 10
D2446 N2446 0 diode
R2447 N2446 N2447 10
D2447 N2447 0 diode
R2448 N2447 N2448 10
D2448 N2448 0 diode
R2449 N2448 N2449 10
D2449 N2449 0 diode
R2450 N2449 N2450 10
D2450 N2450 0 diode
R2451 N2450 N2451 10
D2451 N2451 0 diode
R2452 N2451 N2452 10
D2452 N2452 0 diode
R2453 N2452 N2453 10
D2453 N2453 0 diode
R2454 N2453 N2454 10
D2454 N2454 0 diode
R2455 N2454 N2455 10
D2455 N2455 0 diode
R2456 N2455 N2456 10
D2456 N2456 0 diode
R2457 N2456 N2457 10
D2457 N2457 0 diode
R2458 N2457 N2458 10
D2458 N2458 0 diode
R2459 N2458 N2459 10
D2459 N2459 0 diode
R2460 N2459 N2460 10
D2460 N2460 0 diode
R2461 N2460 N2461 10
D2461 N2461 0 diode
R2462 N2461 N2462 10
D2462 N2462 0 diode
R2463 N2462 N2463 10
D2463 N2463 0 diode
R2464 N2463 N2464 10
D2464 N2464 0 diode
R2465 N2464 N2465 10
D2465 N2465 0 diode
R2466 N2465 N2466 10
D2466 N2466 0 diode
R2467 N2466 N2467 10
D2467 N2467 0 diode
R2468 N2467 N2468 10
D2468 N2468 0 diode
R2469 N2468 N2469 10
D2469 N2469 0 diode
R2470 N2469 N2470 10
D2470 N2470 0 diode
R2471 N2470 N2471 10
D2471 N2471 0 diode
R2472 N2471 N2472 10
D2472 N2472 0 diode
R2473 N2472 N2473 10
D2473 N2473 0 diode
R2474 N2473 N2474 10
D2474 N2474 0 diode
R2475 N2474 N2475 10
D2475 N2475 0 diode
R2476 N2475 N2476 10
D2476 N2476 0 diode
R2477 N2476 N2477 10
D2477 N2477 0 diode
R2478 N2477 N2478 10
D2478 N2478 0 diode
R2479 N2478 N2479 10
D2479 N2479 0 diode
R2480 N2479 N2480 10
D2480 N2480 0 diode
R2481 N2480 N2481 10
D2481 N2481 0 diode
R2482 N2481 N2482 10
D2482 N2482 0 diode
R2483 N2482 N2483 10
D2483 N2483 0 diode
R2484 N2483 N2484 10
D2484 N2484 0 diode
R2485 N2484 N2485 10
D2485 N2485 0 diode
R2486 N2485 N2486 10
D2486 N2486 0 diode
R2487 N2486 N2487 10
D2487 N2487 0 diode
R2488 N2487 N2488 10
D2488 N2488 0 diode
R2489 N2488 N2489 10
D2489 N2489 0 diode
R2490 N2489 N2490 10
D2490 N2490 0 diode
R2491 N2490 N2491 10
D2491 N2491 0 diode
R2492 N2491 N2492 10
D2492 N2492 0 diode
R2493 N2492 N2493 10
D2493 N2493 0 diode
R2494 N2493 N2494 10
D2494 N2494 0 diode
R2495 N2494 N2495 10
D2495 N2495 0 diode
R2496 N2495 N2496 10
D2496 N2496 0 diode
R2497 N2496 N2497 10
D2497 N2497 0 diode
R2498 N2497 N2498 10
D2498 N2498 0 diode
R2499 N2498 N2499 10
D2499 N2499 0 diode
R2500 N2499 N2500 10
D2500 N2500 0 diode
R2501 N2500 N2501 10
D2501 N2501 0 diode
R2502 N2501 N2502 10
D2502 N2502 0 diode
R2503 N2502 N2503 10
D2503 N2503 0 diode
R2504 N2503 N2504 10
D2504 N2504 0 diode
R2505 N2504 N2505 10
D2505 N2505 0 diode
R2506 N2505 N2506 10
D2506 N2506 0 diode
R2507 N2506 N2507 10
D2507 N2507 0 diode
R2508 N2507 N2508 10
D2508 N2508 0 diode
R2509 N2508 N2509 10
D2509 N2509 0 diode
R2510 N2509 N2510 10
D2510 N2510 0 diode
R2511 N2510 N2511 10
D2511 N2511 0 diode
R2512 N2511 N2512 10
D2512 N2512 0 diode
R2513 N2512 N2513 10
D2513 N2513 0 diode
R2514 N2513 N2514 10
D2514 N2514 0 diode
R2515 N2514 N2515 10
D2515 N2515 0 diode
R2516 N2515 N2516 10
D2516 N2516 0 diode
R2517 N2516 N2517 10
D2517 N2517 0 diode
R2518 N2517 N2518 10
D2518 N2518 0 diode
R2519 N2518 N2519 10
D2519 N2519 0 diode
R2520 N2519 N2520 10
D2520 N2520 0 diode
R2521 N2520 N2521 10
D2521 N2521 0 diode
R2522 N2521 N2522 10
D2522 N2522 0 diode
R2523 N2522 N2523 10
D2523 N2523 0 diode
R2524 N2523 N2524 10
D2524 N2524 0 diode
R2525 N2524 N2525 10
D2525 N2525 0 diode
R2526 N2525 N2526 10
D2526 N2526 0 diode
R2527 N2526 N2527 10
D2527 N2527 0 diode
R2528 N2527 N2528 10
D2528 N2528 0 diode
R2529 N2528 N2529 10
D2529 N2529 0 diode
R2530 N2529 N2530 10
D2530 N2530 0 diode
R2531 N2530 N2531 10
D2531 N2531 0 diode
R2532 N2531 N2532 10
D2532 N2532 0 diode
R2533 N2532 N2533 10
D2533 N2533 0 diode
R2534 N2533 N2534 10
D2534 N2534 0 diode
R2535 N2534 N2535 10
D2535 N2535 0 diode
R2536 N2535 N2536 10
D2536 N2536 0 diode
R2537 N2536 N2537 10
D2537 N2537 0 diode
R2538 N2537 N2538 10
D2538 N2538 0 diode
R2539 N2538 N2539 10
D2539 N2539 0 diode
R2540 N2539 N2540 10
D2540 N2540 0 diode
R2541 N2540 N2541 10
D2541 N2541 0 diode
R2542 N2541 N2542 10
D2542 N2542 0 diode
R2543 N2542 N2543 10
D2543 N2543 0 diode
R2544 N2543 N2544 10
D2544 N2544 0 diode
R2545 N2544 N2545 10
D2545 N2545 0 diode
R2546 N2545 N2546 10
D2546 N2546 0 diode
R2547 N2546 N2547 10
D2547 N2547 0 diode
R2548 N2547 N2548 10
D2548 N2548 0 diode
R2549 N2548 N2549 10
D2549 N2549 0 diode
R2550 N2549 N2550 10
D2550 N2550 0 diode
R2551 N2550 N2551 10
D2551 N2551 0 diode
R2552 N2551 N2552 10
D2552 N2552 0 diode
R2553 N2552 N2553 10
D2553 N2553 0 diode
R2554 N2553 N2554 10
D2554 N2554 0 diode
R2555 N2554 N2555 10
D2555 N2555 0 diode
R2556 N2555 N2556 10
D2556 N2556 0 diode
R2557 N2556 N2557 10
D2557 N2557 0 diode
R2558 N2557 N2558 10
D2558 N2558 0 diode
R2559 N2558 N2559 10
D2559 N2559 0 diode
R2560 N2559 N2560 10
D2560 N2560 0 diode
R2561 N2560 N2561 10
D2561 N2561 0 diode
R2562 N2561 N2562 10
D2562 N2562 0 diode
R2563 N2562 N2563 10
D2563 N2563 0 diode
R2564 N2563 N2564 10
D2564 N2564 0 diode
R2565 N2564 N2565 10
D2565 N2565 0 diode
R2566 N2565 N2566 10
D2566 N2566 0 diode
R2567 N2566 N2567 10
D2567 N2567 0 diode
R2568 N2567 N2568 10
D2568 N2568 0 diode
R2569 N2568 N2569 10
D2569 N2569 0 diode
R2570 N2569 N2570 10
D2570 N2570 0 diode
R2571 N2570 N2571 10
D2571 N2571 0 diode
R2572 N2571 N2572 10
D2572 N2572 0 diode
R2573 N2572 N2573 10
D2573 N2573 0 diode
R2574 N2573 N2574 10
D2574 N2574 0 diode
R2575 N2574 N2575 10
D2575 N2575 0 diode
R2576 N2575 N2576 10
D2576 N2576 0 diode
R2577 N2576 N2577 10
D2577 N2577 0 diode
R2578 N2577 N2578 10
D2578 N2578 0 diode
R2579 N2578 N2579 10
D2579 N2579 0 diode
R2580 N2579 N2580 10
D2580 N2580 0 diode
R2581 N2580 N2581 10
D2581 N2581 0 diode
R2582 N2581 N2582 10
D2582 N2582 0 diode
R2583 N2582 N2583 10
D2583 N2583 0 diode
R2584 N2583 N2584 10
D2584 N2584 0 diode
R2585 N2584 N2585 10
D2585 N2585 0 diode
R2586 N2585 N2586 10
D2586 N2586 0 diode
R2587 N2586 N2587 10
D2587 N2587 0 diode
R2588 N2587 N2588 10
D2588 N2588 0 diode
R2589 N2588 N2589 10
D2589 N2589 0 diode
R2590 N2589 N2590 10
D2590 N2590 0 diode
R2591 N2590 N2591 10
D2591 N2591 0 diode
R2592 N2591 N2592 10
D2592 N2592 0 diode
R2593 N2592 N2593 10
D2593 N2593 0 diode
R2594 N2593 N2594 10
D2594 N2594 0 diode
R2595 N2594 N2595 10
D2595 N2595 0 diode
R2596 N2595 N2596 10
D2596 N2596 0 diode
R2597 N2596 N2597 10
D2597 N2597 0 diode
R2598 N2597 N2598 10
D2598 N2598 0 diode
R2599 N2598 N2599 10
D2599 N2599 0 diode
R2600 N2599 N2600 10
D2600 N2600 0 diode
R2601 N2600 N2601 10
D2601 N2601 0 diode
R2602 N2601 N2602 10
D2602 N2602 0 diode
R2603 N2602 N2603 10
D2603 N2603 0 diode
R2604 N2603 N2604 10
D2604 N2604 0 diode
R2605 N2604 N2605 10
D2605 N2605 0 diode
R2606 N2605 N2606 10
D2606 N2606 0 diode
R2607 N2606 N2607 10
D2607 N2607 0 diode
R2608 N2607 N2608 10
D2608 N2608 0 diode
R2609 N2608 N2609 10
D2609 N2609 0 diode
R2610 N2609 N2610 10
D2610 N2610 0 diode
R2611 N2610 N2611 10
D2611 N2611 0 diode
R2612 N2611 N2612 10
D2612 N2612 0 diode
R2613 N2612 N2613 10
D2613 N2613 0 diode
R2614 N2613 N2614 10
D2614 N2614 0 diode
R2615 N2614 N2615 10
D2615 N2615 0 diode
R2616 N2615 N2616 10
D2616 N2616 0 diode
R2617 N2616 N2617 10
D2617 N2617 0 diode
R2618 N2617 N2618 10
D2618 N2618 0 diode
R2619 N2618 N2619 10
D2619 N2619 0 diode
R2620 N2619 N2620 10
D2620 N2620 0 diode
R2621 N2620 N2621 10
D2621 N2621 0 diode
R2622 N2621 N2622 10
D2622 N2622 0 diode
R2623 N2622 N2623 10
D2623 N2623 0 diode
R2624 N2623 N2624 10
D2624 N2624 0 diode
R2625 N2624 N2625 10
D2625 N2625 0 diode
R2626 N2625 N2626 10
D2626 N2626 0 diode
R2627 N2626 N2627 10
D2627 N2627 0 diode
R2628 N2627 N2628 10
D2628 N2628 0 diode
R2629 N2628 N2629 10
D2629 N2629 0 diode
R2630 N2629 N2630 10
D2630 N2630 0 diode
R2631 N2630 N2631 10
D2631 N2631 0 diode
R2632 N2631 N2632 10
D2632 N2632 0 diode
R2633 N2632 N2633 10
D2633 N2633 0 diode
R2634 N2633 N2634 10
D2634 N2634 0 diode
R2635 N2634 N2635 10
D2635 N2635 0 diode
R2636 N2635 N2636 10
D2636 N2636 0 diode
R2637 N2636 N2637 10
D2637 N2637 0 diode
R2638 N2637 N2638 10
D2638 N2638 0 diode
R2639 N2638 N2639 10
D2639 N2639 0 diode
R2640 N2639 N2640 10
D2640 N2640 0 diode
R2641 N2640 N2641 10
D2641 N2641 0 diode
R2642 N2641 N2642 10
D2642 N2642 0 diode
R2643 N2642 N2643 10
D2643 N2643 0 diode
R2644 N2643 N2644 10
D2644 N2644 0 diode
R2645 N2644 N2645 10
D2645 N2645 0 diode
R2646 N2645 N2646 10
D2646 N2646 0 diode
R2647 N2646 N2647 10
D2647 N2647 0 diode
R2648 N2647 N2648 10
D2648 N2648 0 diode
R2649 N2648 N2649 10
D2649 N2649 0 diode
R2650 N2649 N2650 10
D2650 N2650 0 diode
R2651 N2650 N2651 10
D2651 N2651 0 diode
R2652 N2651 N2652 10
D2652 N2652 0 diode
R2653 N2652 N2653 10
D2653 N2653 0 diode
R2654 N2653 N2654 10
D2654 N2654 0 diode
R2655 N2654 N2655 10
D2655 N2655 0 diode
R2656 N2655 N2656 10
D2656 N2656 0 diode
R2657 N2656 N2657 10
D2657 N2657 0 diode
R2658 N2657 N2658 10
D2658 N2658 0 diode
R2659 N2658 N2659 10
D2659 N2659 0 diode
R2660 N2659 N2660 10
D2660 N2660 0 diode
R2661 N2660 N2661 10
D2661 N2661 0 diode
R2662 N2661 N2662 10
D2662 N2662 0 diode
R2663 N2662 N2663 10
D2663 N2663 0 diode
R2664 N2663 N2664 10
D2664 N2664 0 diode
R2665 N2664 N2665 10
D2665 N2665 0 diode
R2666 N2665 N2666 10
D2666 N2666 0 diode
R2667 N2666 N2667 10
D2667 N2667 0 diode
R2668 N2667 N2668 10
D2668 N2668 0 diode
R2669 N2668 N2669 10
D2669 N2669 0 diode
R2670 N2669 N2670 10
D2670 N2670 0 diode
R2671 N2670 N2671 10
D2671 N2671 0 diode
R2672 N2671 N2672 10
D2672 N2672 0 diode
R2673 N2672 N2673 10
D2673 N2673 0 diode
R2674 N2673 N2674 10
D2674 N2674 0 diode
R2675 N2674 N2675 10
D2675 N2675 0 diode
R2676 N2675 N2676 10
D2676 N2676 0 diode
R2677 N2676 N2677 10
D2677 N2677 0 diode
R2678 N2677 N2678 10
D2678 N2678 0 diode
R2679 N2678 N2679 10
D2679 N2679 0 diode
R2680 N2679 N2680 10
D2680 N2680 0 diode
R2681 N2680 N2681 10
D2681 N2681 0 diode
R2682 N2681 N2682 10
D2682 N2682 0 diode
R2683 N2682 N2683 10
D2683 N2683 0 diode
R2684 N2683 N2684 10
D2684 N2684 0 diode
R2685 N2684 N2685 10
D2685 N2685 0 diode
R2686 N2685 N2686 10
D2686 N2686 0 diode
R2687 N2686 N2687 10
D2687 N2687 0 diode
R2688 N2687 N2688 10
D2688 N2688 0 diode
R2689 N2688 N2689 10
D2689 N2689 0 diode
R2690 N2689 N2690 10
D2690 N2690 0 diode
R2691 N2690 N2691 10
D2691 N2691 0 diode
R2692 N2691 N2692 10
D2692 N2692 0 diode
R2693 N2692 N2693 10
D2693 N2693 0 diode
R2694 N2693 N2694 10
D2694 N2694 0 diode
R2695 N2694 N2695 10
D2695 N2695 0 diode
R2696 N2695 N2696 10
D2696 N2696 0 diode
R2697 N2696 N2697 10
D2697 N2697 0 diode
R2698 N2697 N2698 10
D2698 N2698 0 diode
R2699 N2698 N2699 10
D2699 N2699 0 diode
R2700 N2699 N2700 10
D2700 N2700 0 diode
R2701 N2700 N2701 10
D2701 N2701 0 diode
R2702 N2701 N2702 10
D2702 N2702 0 diode
R2703 N2702 N2703 10
D2703 N2703 0 diode
R2704 N2703 N2704 10
D2704 N2704 0 diode
R2705 N2704 N2705 10
D2705 N2705 0 diode
R2706 N2705 N2706 10
D2706 N2706 0 diode
R2707 N2706 N2707 10
D2707 N2707 0 diode
R2708 N2707 N2708 10
D2708 N2708 0 diode
R2709 N2708 N2709 10
D2709 N2709 0 diode
R2710 N2709 N2710 10
D2710 N2710 0 diode
R2711 N2710 N2711 10
D2711 N2711 0 diode
R2712 N2711 N2712 10
D2712 N2712 0 diode
R2713 N2712 N2713 10
D2713 N2713 0 diode
R2714 N2713 N2714 10
D2714 N2714 0 diode
R2715 N2714 N2715 10
D2715 N2715 0 diode
R2716 N2715 N2716 10
D2716 N2716 0 diode
R2717 N2716 N2717 10
D2717 N2717 0 diode
R2718 N2717 N2718 10
D2718 N2718 0 diode
R2719 N2718 N2719 10
D2719 N2719 0 diode
R2720 N2719 N2720 10
D2720 N2720 0 diode
R2721 N2720 N2721 10
D2721 N2721 0 diode
R2722 N2721 N2722 10
D2722 N2722 0 diode
R2723 N2722 N2723 10
D2723 N2723 0 diode
R2724 N2723 N2724 10
D2724 N2724 0 diode
R2725 N2724 N2725 10
D2725 N2725 0 diode
R2726 N2725 N2726 10
D2726 N2726 0 diode
R2727 N2726 N2727 10
D2727 N2727 0 diode
R2728 N2727 N2728 10
D2728 N2728 0 diode
R2729 N2728 N2729 10
D2729 N2729 0 diode
R2730 N2729 N2730 10
D2730 N2730 0 diode
R2731 N2730 N2731 10
D2731 N2731 0 diode
R2732 N2731 N2732 10
D2732 N2732 0 diode
R2733 N2732 N2733 10
D2733 N2733 0 diode
R2734 N2733 N2734 10
D2734 N2734 0 diode
R2735 N2734 N2735 10
D2735 N2735 0 diode
R2736 N2735 N2736 10
D2736 N2736 0 diode
R2737 N2736 N2737 10
D2737 N2737 0 diode
R2738 N2737 N2738 10
D2738 N2738 0 diode
R2739 N2738 N2739 10
D2739 N2739 0 diode
R2740 N2739 N2740 10
D2740 N2740 0 diode
R2741 N2740 N2741 10
D2741 N2741 0 diode
R2742 N2741 N2742 10
D2742 N2742 0 diode
R2743 N2742 N2743 10
D2743 N2743 0 diode
R2744 N2743 N2744 10
D2744 N2744 0 diode
R2745 N2744 N2745 10
D2745 N2745 0 diode
R2746 N2745 N2746 10
D2746 N2746 0 diode
R2747 N2746 N2747 10
D2747 N2747 0 diode
R2748 N2747 N2748 10
D2748 N2748 0 diode
R2749 N2748 N2749 10
D2749 N2749 0 diode
R2750 N2749 N2750 10
D2750 N2750 0 diode
R2751 N2750 N2751 10
D2751 N2751 0 diode
R2752 N2751 N2752 10
D2752 N2752 0 diode
R2753 N2752 N2753 10
D2753 N2753 0 diode
R2754 N2753 N2754 10
D2754 N2754 0 diode
R2755 N2754 N2755 10
D2755 N2755 0 diode
R2756 N2755 N2756 10
D2756 N2756 0 diode
R2757 N2756 N2757 10
D2757 N2757 0 diode
R2758 N2757 N2758 10
D2758 N2758 0 diode
R2759 N2758 N2759 10
D2759 N2759 0 diode
R2760 N2759 N2760 10
D2760 N2760 0 diode
R2761 N2760 N2761 10
D2761 N2761 0 diode
R2762 N2761 N2762 10
D2762 N2762 0 diode
R2763 N2762 N2763 10
D2763 N2763 0 diode
R2764 N2763 N2764 10
D2764 N2764 0 diode
R2765 N2764 N2765 10
D2765 N2765 0 diode
R2766 N2765 N2766 10
D2766 N2766 0 diode
R2767 N2766 N2767 10
D2767 N2767 0 diode
R2768 N2767 N2768 10
D2768 N2768 0 diode
R2769 N2768 N2769 10
D2769 N2769 0 diode
R2770 N2769 N2770 10
D2770 N2770 0 diode
R2771 N2770 N2771 10
D2771 N2771 0 diode
R2772 N2771 N2772 10
D2772 N2772 0 diode
R2773 N2772 N2773 10
D2773 N2773 0 diode
R2774 N2773 N2774 10
D2774 N2774 0 diode
R2775 N2774 N2775 10
D2775 N2775 0 diode
R2776 N2775 N2776 10
D2776 N2776 0 diode
R2777 N2776 N2777 10
D2777 N2777 0 diode
R2778 N2777 N2778 10
D2778 N2778 0 diode
R2779 N2778 N2779 10
D2779 N2779 0 diode
R2780 N2779 N2780 10
D2780 N2780 0 diode
R2781 N2780 N2781 10
D2781 N2781 0 diode
R2782 N2781 N2782 10
D2782 N2782 0 diode
R2783 N2782 N2783 10
D2783 N2783 0 diode
R2784 N2783 N2784 10
D2784 N2784 0 diode
R2785 N2784 N2785 10
D2785 N2785 0 diode
R2786 N2785 N2786 10
D2786 N2786 0 diode
R2787 N2786 N2787 10
D2787 N2787 0 diode
R2788 N2787 N2788 10
D2788 N2788 0 diode
R2789 N2788 N2789 10
D2789 N2789 0 diode
R2790 N2789 N2790 10
D2790 N2790 0 diode
R2791 N2790 N2791 10
D2791 N2791 0 diode
R2792 N2791 N2792 10
D2792 N2792 0 diode
R2793 N2792 N2793 10
D2793 N2793 0 diode
R2794 N2793 N2794 10
D2794 N2794 0 diode
R2795 N2794 N2795 10
D2795 N2795 0 diode
R2796 N2795 N2796 10
D2796 N2796 0 diode
R2797 N2796 N2797 10
D2797 N2797 0 diode
R2798 N2797 N2798 10
D2798 N2798 0 diode
R2799 N2798 N2799 10
D2799 N2799 0 diode
R2800 N2799 N2800 10
D2800 N2800 0 diode
R2801 N2800 N2801 10
D2801 N2801 0 diode
R2802 N2801 N2802 10
D2802 N2802 0 diode
R2803 N2802 N2803 10
D2803 N2803 0 diode
R2804 N2803 N2804 10
D2804 N2804 0 diode
R2805 N2804 N2805 10
D2805 N2805 0 diode
R2806 N2805 N2806 10
D2806 N2806 0 diode
R2807 N2806 N2807 10
D2807 N2807 0 diode
R2808 N2807 N2808 10
D2808 N2808 0 diode
R2809 N2808 N2809 10
D2809 N2809 0 diode
R2810 N2809 N2810 10
D2810 N2810 0 diode
R2811 N2810 N2811 10
D2811 N2811 0 diode
R2812 N2811 N2812 10
D2812 N2812 0 diode
R2813 N2812 N2813 10
D2813 N2813 0 diode
R2814 N2813 N2814 10
D2814 N2814 0 diode
R2815 N2814 N2815 10
D2815 N2815 0 diode
R2816 N2815 N2816 10
D2816 N2816 0 diode
R2817 N2816 N2817 10
D2817 N2817 0 diode
R2818 N2817 N2818 10
D2818 N2818 0 diode
R2819 N2818 N2819 10
D2819 N2819 0 diode
R2820 N2819 N2820 10
D2820 N2820 0 diode
R2821 N2820 N2821 10
D2821 N2821 0 diode
R2822 N2821 N2822 10
D2822 N2822 0 diode
R2823 N2822 N2823 10
D2823 N2823 0 diode
R2824 N2823 N2824 10
D2824 N2824 0 diode
R2825 N2824 N2825 10
D2825 N2825 0 diode
R2826 N2825 N2826 10
D2826 N2826 0 diode
R2827 N2826 N2827 10
D2827 N2827 0 diode
R2828 N2827 N2828 10
D2828 N2828 0 diode
R2829 N2828 N2829 10
D2829 N2829 0 diode
R2830 N2829 N2830 10
D2830 N2830 0 diode
R2831 N2830 N2831 10
D2831 N2831 0 diode
R2832 N2831 N2832 10
D2832 N2832 0 diode
R2833 N2832 N2833 10
D2833 N2833 0 diode
R2834 N2833 N2834 10
D2834 N2834 0 diode
R2835 N2834 N2835 10
D2835 N2835 0 diode
R2836 N2835 N2836 10
D2836 N2836 0 diode
R2837 N2836 N2837 10
D2837 N2837 0 diode
R2838 N2837 N2838 10
D2838 N2838 0 diode
R2839 N2838 N2839 10
D2839 N2839 0 diode
R2840 N2839 N2840 10
D2840 N2840 0 diode
R2841 N2840 N2841 10
D2841 N2841 0 diode
R2842 N2841 N2842 10
D2842 N2842 0 diode
R2843 N2842 N2843 10
D2843 N2843 0 diode
R2844 N2843 N2844 10
D2844 N2844 0 diode
R2845 N2844 N2845 10
D2845 N2845 0 diode
R2846 N2845 N2846 10
D2846 N2846 0 diode
R2847 N2846 N2847 10
D2847 N2847 0 diode
R2848 N2847 N2848 10
D2848 N2848 0 diode
R2849 N2848 N2849 10
D2849 N2849 0 diode
R2850 N2849 N2850 10
D2850 N2850 0 diode
R2851 N2850 N2851 10
D2851 N2851 0 diode
R2852 N2851 N2852 10
D2852 N2852 0 diode
R2853 N2852 N2853 10
D2853 N2853 0 diode
R2854 N2853 N2854 10
D2854 N2854 0 diode
R2855 N2854 N2855 10
D2855 N2855 0 diode
R2856 N2855 N2856 10
D2856 N2856 0 diode
R2857 N2856 N2857 10
D2857 N2857 0 diode
R2858 N2857 N2858 10
D2858 N2858 0 diode
R2859 N2858 N2859 10
D2859 N2859 0 diode
R2860 N2859 N2860 10
D2860 N2860 0 diode
R2861 N2860 N2861 10
D2861 N2861 0 diode
R2862 N2861 N2862 10
D2862 N2862 0 diode
R2863 N2862 N2863 10
D2863 N2863 0 diode
R2864 N2863 N2864 10
D2864 N2864 0 diode
R2865 N2864 N2865 10
D2865 N2865 0 diode
R2866 N2865 N2866 10
D2866 N2866 0 diode
R2867 N2866 N2867 10
D2867 N2867 0 diode
R2868 N2867 N2868 10
D2868 N2868 0 diode
R2869 N2868 N2869 10
D2869 N2869 0 diode
R2870 N2869 N2870 10
D2870 N2870 0 diode
R2871 N2870 N2871 10
D2871 N2871 0 diode
R2872 N2871 N2872 10
D2872 N2872 0 diode
R2873 N2872 N2873 10
D2873 N2873 0 diode
R2874 N2873 N2874 10
D2874 N2874 0 diode
R2875 N2874 N2875 10
D2875 N2875 0 diode
R2876 N2875 N2876 10
D2876 N2876 0 diode
R2877 N2876 N2877 10
D2877 N2877 0 diode
R2878 N2877 N2878 10
D2878 N2878 0 diode
R2879 N2878 N2879 10
D2879 N2879 0 diode
R2880 N2879 N2880 10
D2880 N2880 0 diode
R2881 N2880 N2881 10
D2881 N2881 0 diode
R2882 N2881 N2882 10
D2882 N2882 0 diode
R2883 N2882 N2883 10
D2883 N2883 0 diode
R2884 N2883 N2884 10
D2884 N2884 0 diode
R2885 N2884 N2885 10
D2885 N2885 0 diode
R2886 N2885 N2886 10
D2886 N2886 0 diode
R2887 N2886 N2887 10
D2887 N2887 0 diode
R2888 N2887 N2888 10
D2888 N2888 0 diode
R2889 N2888 N2889 10
D2889 N2889 0 diode
R2890 N2889 N2890 10
D2890 N2890 0 diode
R2891 N2890 N2891 10
D2891 N2891 0 diode
R2892 N2891 N2892 10
D2892 N2892 0 diode
R2893 N2892 N2893 10
D2893 N2893 0 diode
R2894 N2893 N2894 10
D2894 N2894 0 diode
R2895 N2894 N2895 10
D2895 N2895 0 diode
R2896 N2895 N2896 10
D2896 N2896 0 diode
R2897 N2896 N2897 10
D2897 N2897 0 diode
R2898 N2897 N2898 10
D2898 N2898 0 diode
R2899 N2898 N2899 10
D2899 N2899 0 diode
R2900 N2899 N2900 10
D2900 N2900 0 diode
R2901 N2900 N2901 10
D2901 N2901 0 diode
R2902 N2901 N2902 10
D2902 N2902 0 diode
R2903 N2902 N2903 10
D2903 N2903 0 diode
R2904 N2903 N2904 10
D2904 N2904 0 diode
R2905 N2904 N2905 10
D2905 N2905 0 diode
R2906 N2905 N2906 10
D2906 N2906 0 diode
R2907 N2906 N2907 10
D2907 N2907 0 diode
R2908 N2907 N2908 10
D2908 N2908 0 diode
R2909 N2908 N2909 10
D2909 N2909 0 diode
R2910 N2909 N2910 10
D2910 N2910 0 diode
R2911 N2910 N2911 10
D2911 N2911 0 diode
R2912 N2911 N2912 10
D2912 N2912 0 diode
R2913 N2912 N2913 10
D2913 N2913 0 diode
R2914 N2913 N2914 10
D2914 N2914 0 diode
R2915 N2914 N2915 10
D2915 N2915 0 diode
R2916 N2915 N2916 10
D2916 N2916 0 diode
R2917 N2916 N2917 10
D2917 N2917 0 diode
R2918 N2917 N2918 10
D2918 N2918 0 diode
R2919 N2918 N2919 10
D2919 N2919 0 diode
R2920 N2919 N2920 10
D2920 N2920 0 diode
R2921 N2920 N2921 10
D2921 N2921 0 diode
R2922 N2921 N2922 10
D2922 N2922 0 diode
R2923 N2922 N2923 10
D2923 N2923 0 diode
R2924 N2923 N2924 10
D2924 N2924 0 diode
R2925 N2924 N2925 10
D2925 N2925 0 diode
R2926 N2925 N2926 10
D2926 N2926 0 diode
R2927 N2926 N2927 10
D2927 N2927 0 diode
R2928 N2927 N2928 10
D2928 N2928 0 diode
R2929 N2928 N2929 10
D2929 N2929 0 diode
R2930 N2929 N2930 10
D2930 N2930 0 diode
R2931 N2930 N2931 10
D2931 N2931 0 diode
R2932 N2931 N2932 10
D2932 N2932 0 diode
R2933 N2932 N2933 10
D2933 N2933 0 diode
R2934 N2933 N2934 10
D2934 N2934 0 diode
R2935 N2934 N2935 10
D2935 N2935 0 diode
R2936 N2935 N2936 10
D2936 N2936 0 diode
R2937 N2936 N2937 10
D2937 N2937 0 diode
R2938 N2937 N2938 10
D2938 N2938 0 diode
R2939 N2938 N2939 10
D2939 N2939 0 diode
R2940 N2939 N2940 10
D2940 N2940 0 diode
R2941 N2940 N2941 10
D2941 N2941 0 diode
R2942 N2941 N2942 10
D2942 N2942 0 diode
R2943 N2942 N2943 10
D2943 N2943 0 diode
R2944 N2943 N2944 10
D2944 N2944 0 diode
R2945 N2944 N2945 10
D2945 N2945 0 diode
R2946 N2945 N2946 10
D2946 N2946 0 diode
R2947 N2946 N2947 10
D2947 N2947 0 diode
R2948 N2947 N2948 10
D2948 N2948 0 diode
R2949 N2948 N2949 10
D2949 N2949 0 diode
R2950 N2949 N2950 10
D2950 N2950 0 diode
R2951 N2950 N2951 10
D2951 N2951 0 diode
R2952 N2951 N2952 10
D2952 N2952 0 diode
R2953 N2952 N2953 10
D2953 N2953 0 diode
R2954 N2953 N2954 10
D2954 N2954 0 diode
R2955 N2954 N2955 10
D2955 N2955 0 diode
R2956 N2955 N2956 10
D2956 N2956 0 diode
R2957 N2956 N2957 10
D2957 N2957 0 diode
R2958 N2957 N2958 10
D2958 N2958 0 diode
R2959 N2958 N2959 10
D2959 N2959 0 diode
R2960 N2959 N2960 10
D2960 N2960 0 diode
R2961 N2960 N2961 10
D2961 N2961 0 diode
R2962 N2961 N2962 10
D2962 N2962 0 diode
R2963 N2962 N2963 10
D2963 N2963 0 diode
R2964 N2963 N2964 10
D2964 N2964 0 diode
R2965 N2964 N2965 10
D2965 N2965 0 diode
R2966 N2965 N2966 10
D2966 N2966 0 diode
R2967 N2966 N2967 10
D2967 N2967 0 diode
R2968 N2967 N2968 10
D2968 N2968 0 diode
R2969 N2968 N2969 10
D2969 N2969 0 diode
R2970 N2969 N2970 10
D2970 N2970 0 diode
R2971 N2970 N2971 10
D2971 N2971 0 diode
R2972 N2971 N2972 10
D2972 N2972 0 diode
R2973 N2972 N2973 10
D2973 N2973 0 diode
R2974 N2973 N2974 10
D2974 N2974 0 diode
R2975 N2974 N2975 10
D2975 N2975 0 diode
R2976 N2975 N2976 10
D2976 N2976 0 diode
R2977 N2976 N2977 10
D2977 N2977 0 diode
R2978 N2977 N2978 10
D2978 N2978 0 diode
R2979 N2978 N2979 10
D2979 N2979 0 diode
R2980 N2979 N2980 10
D2980 N2980 0 diode
R2981 N2980 N2981 10
D2981 N2981 0 diode
R2982 N2981 N2982 10
D2982 N2982 0 diode
R2983 N2982 N2983 10
D2983 N2983 0 diode
R2984 N2983 N2984 10
D2984 N2984 0 diode
R2985 N2984 N2985 10
D2985 N2985 0 diode
R2986 N2985 N2986 10
D2986 N2986 0 diode
R2987 N2986 N2987 10
D2987 N2987 0 diode
R2988 N2987 N2988 10
D2988 N2988 0 diode
R2989 N2988 N2989 10
D2989 N2989 0 diode
R2990 N2989 N2990 10
D2990 N2990 0 diode
R2991 N2990 N2991 10
D2991 N2991 0 diode
R2992 N2991 N2992 10
D2992 N2992 0 diode
R2993 N2992 N2993 10
D2993 N2993 0 diode
R2994 N2993 N2994 10
D2994 N2994 0 diode
R2995 N2994 N2995 10
D2995 N2995 0 diode
R2996 N2995 N2996 10
D2996 N2996 0 diode
R2997 N2996 N2997 10
D2997 N2997 0 diode
R2998 N2997 N2998 10
D2998 N2998 0 diode
R2999 N2998 N2999 10
D2999 N2999 0 diode
R3000 N2999 N3000 10
D3000 N3000 0 diode
R3001 N3000 N3001 10
D3001 N3001 0 diode
R3002 N3001 N3002 10
D3002 N3002 0 diode
R3003 N3002 N3003 10
D3003 N3003 0 diode
R3004 N3003 N3004 10
D3004 N3004 0 diode
R3005 N3004 N3005 10
D3005 N3005 0 diode
R3006 N3005 N3006 10
D3006 N3006 0 diode
R3007 N3006 N3007 10
D3007 N3007 0 diode
R3008 N3007 N3008 10
D3008 N3008 0 diode
R3009 N3008 N3009 10
D3009 N3009 0 diode
R3010 N3009 N3010 10
D3010 N3010 0 diode
R3011 N3010 N3011 10
D3011 N3011 0 diode
R3012 N3011 N3012 10
D3012 N3012 0 diode
R3013 N3012 N3013 10
D3013 N3013 0 diode
R3014 N3013 N3014 10
D3014 N3014 0 diode
R3015 N3014 N3015 10
D3015 N3015 0 diode
R3016 N3015 N3016 10
D3016 N3016 0 diode
R3017 N3016 N3017 10
D3017 N3017 0 diode
R3018 N3017 N3018 10
D3018 N3018 0 diode
R3019 N3018 N3019 10
D3019 N3019 0 diode
R3020 N3019 N3020 10
D3020 N3020 0 diode
R3021 N3020 N3021 10
D3021 N3021 0 diode
R3022 N3021 N3022 10
D3022 N3022 0 diode
R3023 N3022 N3023 10
D3023 N3023 0 diode
R3024 N3023 N3024 10
D3024 N3024 0 diode
R3025 N3024 N3025 10
D3025 N3025 0 diode
R3026 N3025 N3026 10
D3026 N3026 0 diode
R3027 N3026 N3027 10
D3027 N3027 0 diode
R3028 N3027 N3028 10
D3028 N3028 0 diode
R3029 N3028 N3029 10
D3029 N3029 0 diode
R3030 N3029 N3030 10
D3030 N3030 0 diode
R3031 N3030 N3031 10
D3031 N3031 0 diode
R3032 N3031 N3032 10
D3032 N3032 0 diode
R3033 N3032 N3033 10
D3033 N3033 0 diode
R3034 N3033 N3034 10
D3034 N3034 0 diode
R3035 N3034 N3035 10
D3035 N3035 0 diode
R3036 N3035 N3036 10
D3036 N3036 0 diode
R3037 N3036 N3037 10
D3037 N3037 0 diode
R3038 N3037 N3038 10
D3038 N3038 0 diode
R3039 N3038 N3039 10
D3039 N3039 0 diode
R3040 N3039 N3040 10
D3040 N3040 0 diode
R3041 N3040 N3041 10
D3041 N3041 0 diode
R3042 N3041 N3042 10
D3042 N3042 0 diode
R3043 N3042 N3043 10
D3043 N3043 0 diode
R3044 N3043 N3044 10
D3044 N3044 0 diode
R3045 N3044 N3045 10
D3045 N3045 0 diode
R3046 N3045 N3046 10
D3046 N3046 0 diode
R3047 N3046 N3047 10
D3047 N3047 0 diode
R3048 N3047 N3048 10
D3048 N3048 0 diode
R3049 N3048 N3049 10
D3049 N3049 0 diode
R3050 N3049 N3050 10
D3050 N3050 0 diode
R3051 N3050 N3051 10
D3051 N3051 0 diode
R3052 N3051 N3052 10
D3052 N3052 0 diode
R3053 N3052 N3053 10
D3053 N3053 0 diode
R3054 N3053 N3054 10
D3054 N3054 0 diode
R3055 N3054 N3055 10
D3055 N3055 0 diode
R3056 N3055 N3056 10
D3056 N3056 0 diode
R3057 N3056 N3057 10
D3057 N3057 0 diode
R3058 N3057 N3058 10
D3058 N3058 0 diode
R3059 N3058 N3059 10
D3059 N3059 0 diode
R3060 N3059 N3060 10
D3060 N3060 0 diode
R3061 N3060 N3061 10
D3061 N3061 0 diode
R3062 N3061 N3062 10
D3062 N3062 0 diode
R3063 N3062 N3063 10
D3063 N3063 0 diode
R3064 N3063 N3064 10
D3064 N3064 0 diode
R3065 N3064 N3065 10
D3065 N3065 0 diode
R3066 N3065 N3066 10
D3066 N3066 0 diode
R3067 N3066 N3067 10
D3067 N3067 0 diode
R3068 N3067 N3068 10
D3068 N3068 0 diode
R3069 N3068 N3069 10
D3069 N3069 0 diode
R3070 N3069 N3070 10
D3070 N3070 0 diode
R3071 N3070 N3071 10
D3071 N3071 0 diode
R3072 N3071 N3072 10
D3072 N3072 0 diode
R3073 N3072 N3073 10
D3073 N3073 0 diode
R3074 N3073 N3074 10
D3074 N3074 0 diode
R3075 N3074 N3075 10
D3075 N3075 0 diode
R3076 N3075 N3076 10
D3076 N3076 0 diode
R3077 N3076 N3077 10
D3077 N3077 0 diode
R3078 N3077 N3078 10
D3078 N3078 0 diode
R3079 N3078 N3079 10
D3079 N3079 0 diode
R3080 N3079 N3080 10
D3080 N3080 0 diode
R3081 N3080 N3081 10
D3081 N3081 0 diode
R3082 N3081 N3082 10
D3082 N3082 0 diode
R3083 N3082 N3083 10
D3083 N3083 0 diode
R3084 N3083 N3084 10
D3084 N3084 0 diode
R3085 N3084 N3085 10
D3085 N3085 0 diode
R3086 N3085 N3086 10
D3086 N3086 0 diode
R3087 N3086 N3087 10
D3087 N3087 0 diode
R3088 N3087 N3088 10
D3088 N3088 0 diode
R3089 N3088 N3089 10
D3089 N3089 0 diode
R3090 N3089 N3090 10
D3090 N3090 0 diode
R3091 N3090 N3091 10
D3091 N3091 0 diode
R3092 N3091 N3092 10
D3092 N3092 0 diode
R3093 N3092 N3093 10
D3093 N3093 0 diode
R3094 N3093 N3094 10
D3094 N3094 0 diode
R3095 N3094 N3095 10
D3095 N3095 0 diode
R3096 N3095 N3096 10
D3096 N3096 0 diode
R3097 N3096 N3097 10
D3097 N3097 0 diode
R3098 N3097 N3098 10
D3098 N3098 0 diode
R3099 N3098 N3099 10
D3099 N3099 0 diode
R3100 N3099 N3100 10
D3100 N3100 0 diode
R3101 N3100 N3101 10
D3101 N3101 0 diode
R3102 N3101 N3102 10
D3102 N3102 0 diode
R3103 N3102 N3103 10
D3103 N3103 0 diode
R3104 N3103 N3104 10
D3104 N3104 0 diode
R3105 N3104 N3105 10
D3105 N3105 0 diode
R3106 N3105 N3106 10
D3106 N3106 0 diode
R3107 N3106 N3107 10
D3107 N3107 0 diode
R3108 N3107 N3108 10
D3108 N3108 0 diode
R3109 N3108 N3109 10
D3109 N3109 0 diode
R3110 N3109 N3110 10
D3110 N3110 0 diode
R3111 N3110 N3111 10
D3111 N3111 0 diode
R3112 N3111 N3112 10
D3112 N3112 0 diode
R3113 N3112 N3113 10
D3113 N3113 0 diode
R3114 N3113 N3114 10
D3114 N3114 0 diode
R3115 N3114 N3115 10
D3115 N3115 0 diode
R3116 N3115 N3116 10
D3116 N3116 0 diode
R3117 N3116 N3117 10
D3117 N3117 0 diode
R3118 N3117 N3118 10
D3118 N3118 0 diode
R3119 N3118 N3119 10
D3119 N3119 0 diode
R3120 N3119 N3120 10
D3120 N3120 0 diode
R3121 N3120 N3121 10
D3121 N3121 0 diode
R3122 N3121 N3122 10
D3122 N3122 0 diode
R3123 N3122 N3123 10
D3123 N3123 0 diode
R3124 N3123 N3124 10
D3124 N3124 0 diode
R3125 N3124 N3125 10
D3125 N3125 0 diode
R3126 N3125 N3126 10
D3126 N3126 0 diode
R3127 N3126 N3127 10
D3127 N3127 0 diode
R3128 N3127 N3128 10
D3128 N3128 0 diode
R3129 N3128 N3129 10
D3129 N3129 0 diode
R3130 N3129 N3130 10
D3130 N3130 0 diode
R3131 N3130 N3131 10
D3131 N3131 0 diode
R3132 N3131 N3132 10
D3132 N3132 0 diode
R3133 N3132 N3133 10
D3133 N3133 0 diode
R3134 N3133 N3134 10
D3134 N3134 0 diode
R3135 N3134 N3135 10
D3135 N3135 0 diode
R3136 N3135 N3136 10
D3136 N3136 0 diode
R3137 N3136 N3137 10
D3137 N3137 0 diode
R3138 N3137 N3138 10
D3138 N3138 0 diode
R3139 N3138 N3139 10
D3139 N3139 0 diode
R3140 N3139 N3140 10
D3140 N3140 0 diode
R3141 N3140 N3141 10
D3141 N3141 0 diode
R3142 N3141 N3142 10
D3142 N3142 0 diode
R3143 N3142 N3143 10
D3143 N3143 0 diode
R3144 N3143 N3144 10
D3144 N3144 0 diode
R3145 N3144 N3145 10
D3145 N3145 0 diode
R3146 N3145 N3146 10
D3146 N3146 0 diode
R3147 N3146 N3147 10
D3147 N3147 0 diode
R3148 N3147 N3148 10
D3148 N3148 0 diode
R3149 N3148 N3149 10
D3149 N3149 0 diode
R3150 N3149 N3150 10
D3150 N3150 0 diode
R3151 N3150 N3151 10
D3151 N3151 0 diode
R3152 N3151 N3152 10
D3152 N3152 0 diode
R3153 N3152 N3153 10
D3153 N3153 0 diode
R3154 N3153 N3154 10
D3154 N3154 0 diode
R3155 N3154 N3155 10
D3155 N3155 0 diode
R3156 N3155 N3156 10
D3156 N3156 0 diode
R3157 N3156 N3157 10
D3157 N3157 0 diode
R3158 N3157 N3158 10
D3158 N3158 0 diode
R3159 N3158 N3159 10
D3159 N3159 0 diode
R3160 N3159 N3160 10
D3160 N3160 0 diode
R3161 N3160 N3161 10
D3161 N3161 0 diode
R3162 N3161 N3162 10
D3162 N3162 0 diode
R3163 N3162 N3163 10
D3163 N3163 0 diode
R3164 N3163 N3164 10
D3164 N3164 0 diode
R3165 N3164 N3165 10
D3165 N3165 0 diode
R3166 N3165 N3166 10
D3166 N3166 0 diode
R3167 N3166 N3167 10
D3167 N3167 0 diode
R3168 N3167 N3168 10
D3168 N3168 0 diode
R3169 N3168 N3169 10
D3169 N3169 0 diode
R3170 N3169 N3170 10
D3170 N3170 0 diode
R3171 N3170 N3171 10
D3171 N3171 0 diode
R3172 N3171 N3172 10
D3172 N3172 0 diode
R3173 N3172 N3173 10
D3173 N3173 0 diode
R3174 N3173 N3174 10
D3174 N3174 0 diode
R3175 N3174 N3175 10
D3175 N3175 0 diode
R3176 N3175 N3176 10
D3176 N3176 0 diode
R3177 N3176 N3177 10
D3177 N3177 0 diode
R3178 N3177 N3178 10
D3178 N3178 0 diode
R3179 N3178 N3179 10
D3179 N3179 0 diode
R3180 N3179 N3180 10
D3180 N3180 0 diode
R3181 N3180 N3181 10
D3181 N3181 0 diode
R3182 N3181 N3182 10
D3182 N3182 0 diode
R3183 N3182 N3183 10
D3183 N3183 0 diode
R3184 N3183 N3184 10
D3184 N3184 0 diode
R3185 N3184 N3185 10
D3185 N3185 0 diode
R3186 N3185 N3186 10
D3186 N3186 0 diode
R3187 N3186 N3187 10
D3187 N3187 0 diode
R3188 N3187 N3188 10
D3188 N3188 0 diode
R3189 N3188 N3189 10
D3189 N3189 0 diode
R3190 N3189 N3190 10
D3190 N3190 0 diode
R3191 N3190 N3191 10
D3191 N3191 0 diode
R3192 N3191 N3192 10
D3192 N3192 0 diode
R3193 N3192 N3193 10
D3193 N3193 0 diode
R3194 N3193 N3194 10
D3194 N3194 0 diode
R3195 N3194 N3195 10
D3195 N3195 0 diode
R3196 N3195 N3196 10
D3196 N3196 0 diode
R3197 N3196 N3197 10
D3197 N3197 0 diode
R3198 N3197 N3198 10
D3198 N3198 0 diode
R3199 N3198 N3199 10
D3199 N3199 0 diode
R3200 N3199 N3200 10
D3200 N3200 0 diode
R3201 N3200 N3201 10
D3201 N3201 0 diode
R3202 N3201 N3202 10
D3202 N3202 0 diode
R3203 N3202 N3203 10
D3203 N3203 0 diode
R3204 N3203 N3204 10
D3204 N3204 0 diode
R3205 N3204 N3205 10
D3205 N3205 0 diode
R3206 N3205 N3206 10
D3206 N3206 0 diode
R3207 N3206 N3207 10
D3207 N3207 0 diode
R3208 N3207 N3208 10
D3208 N3208 0 diode
R3209 N3208 N3209 10
D3209 N3209 0 diode
R3210 N3209 N3210 10
D3210 N3210 0 diode
R3211 N3210 N3211 10
D3211 N3211 0 diode
R3212 N3211 N3212 10
D3212 N3212 0 diode
R3213 N3212 N3213 10
D3213 N3213 0 diode
R3214 N3213 N3214 10
D3214 N3214 0 diode
R3215 N3214 N3215 10
D3215 N3215 0 diode
R3216 N3215 N3216 10
D3216 N3216 0 diode
R3217 N3216 N3217 10
D3217 N3217 0 diode
R3218 N3217 N3218 10
D3218 N3218 0 diode
R3219 N3218 N3219 10
D3219 N3219 0 diode
R3220 N3219 N3220 10
D3220 N3220 0 diode
R3221 N3220 N3221 10
D3221 N3221 0 diode
R3222 N3221 N3222 10
D3222 N3222 0 diode
R3223 N3222 N3223 10
D3223 N3223 0 diode
R3224 N3223 N3224 10
D3224 N3224 0 diode
R3225 N3224 N3225 10
D3225 N3225 0 diode
R3226 N3225 N3226 10
D3226 N3226 0 diode
R3227 N3226 N3227 10
D3227 N3227 0 diode
R3228 N3227 N3228 10
D3228 N3228 0 diode
R3229 N3228 N3229 10
D3229 N3229 0 diode
R3230 N3229 N3230 10
D3230 N3230 0 diode
R3231 N3230 N3231 10
D3231 N3231 0 diode
R3232 N3231 N3232 10
D3232 N3232 0 diode
R3233 N3232 N3233 10
D3233 N3233 0 diode
R3234 N3233 N3234 10
D3234 N3234 0 diode
R3235 N3234 N3235 10
D3235 N3235 0 diode
R3236 N3235 N3236 10
D3236 N3236 0 diode
R3237 N3236 N3237 10
D3237 N3237 0 diode
R3238 N3237 N3238 10
D3238 N3238 0 diode
R3239 N3238 N3239 10
D3239 N3239 0 diode
R3240 N3239 N3240 10
D3240 N3240 0 diode
R3241 N3240 N3241 10
D3241 N3241 0 diode
R3242 N3241 N3242 10
D3242 N3242 0 diode
R3243 N3242 N3243 10
D3243 N3243 0 diode
R3244 N3243 N3244 10
D3244 N3244 0 diode
R3245 N3244 N3245 10
D3245 N3245 0 diode
R3246 N3245 N3246 10
D3246 N3246 0 diode
R3247 N3246 N3247 10
D3247 N3247 0 diode
R3248 N3247 N3248 10
D3248 N3248 0 diode
R3249 N3248 N3249 10
D3249 N3249 0 diode
R3250 N3249 N3250 10
D3250 N3250 0 diode
R3251 N3250 N3251 10
D3251 N3251 0 diode
R3252 N3251 N3252 10
D3252 N3252 0 diode
R3253 N3252 N3253 10
D3253 N3253 0 diode
R3254 N3253 N3254 10
D3254 N3254 0 diode
R3255 N3254 N3255 10
D3255 N3255 0 diode
R3256 N3255 N3256 10
D3256 N3256 0 diode
R3257 N3256 N3257 10
D3257 N3257 0 diode
R3258 N3257 N3258 10
D3258 N3258 0 diode
R3259 N3258 N3259 10
D3259 N3259 0 diode
R3260 N3259 N3260 10
D3260 N3260 0 diode
R3261 N3260 N3261 10
D3261 N3261 0 diode
R3262 N3261 N3262 10
D3262 N3262 0 diode
R3263 N3262 N3263 10
D3263 N3263 0 diode
R3264 N3263 N3264 10
D3264 N3264 0 diode
R3265 N3264 N3265 10
D3265 N3265 0 diode
R3266 N3265 N3266 10
D3266 N3266 0 diode
R3267 N3266 N3267 10
D3267 N3267 0 diode
R3268 N3267 N3268 10
D3268 N3268 0 diode
R3269 N3268 N3269 10
D3269 N3269 0 diode
R3270 N3269 N3270 10
D3270 N3270 0 diode
R3271 N3270 N3271 10
D3271 N3271 0 diode
R3272 N3271 N3272 10
D3272 N3272 0 diode
R3273 N3272 N3273 10
D3273 N3273 0 diode
R3274 N3273 N3274 10
D3274 N3274 0 diode
R3275 N3274 N3275 10
D3275 N3275 0 diode
R3276 N3275 N3276 10
D3276 N3276 0 diode
R3277 N3276 N3277 10
D3277 N3277 0 diode
R3278 N3277 N3278 10
D3278 N3278 0 diode
R3279 N3278 N3279 10
D3279 N3279 0 diode
R3280 N3279 N3280 10
D3280 N3280 0 diode
R3281 N3280 N3281 10
D3281 N3281 0 diode
R3282 N3281 N3282 10
D3282 N3282 0 diode
R3283 N3282 N3283 10
D3283 N3283 0 diode
R3284 N3283 N3284 10
D3284 N3284 0 diode
R3285 N3284 N3285 10
D3285 N3285 0 diode
R3286 N3285 N3286 10
D3286 N3286 0 diode
R3287 N3286 N3287 10
D3287 N3287 0 diode
R3288 N3287 N3288 10
D3288 N3288 0 diode
R3289 N3288 N3289 10
D3289 N3289 0 diode
R3290 N3289 N3290 10
D3290 N3290 0 diode
R3291 N3290 N3291 10
D3291 N3291 0 diode
R3292 N3291 N3292 10
D3292 N3292 0 diode
R3293 N3292 N3293 10
D3293 N3293 0 diode
R3294 N3293 N3294 10
D3294 N3294 0 diode
R3295 N3294 N3295 10
D3295 N3295 0 diode
R3296 N3295 N3296 10
D3296 N3296 0 diode
R3297 N3296 N3297 10
D3297 N3297 0 diode
R3298 N3297 N3298 10
D3298 N3298 0 diode
R3299 N3298 N3299 10
D3299 N3299 0 diode
R3300 N3299 N3300 10
D3300 N3300 0 diode
R3301 N3300 N3301 10
D3301 N3301 0 diode
R3302 N3301 N3302 10
D3302 N3302 0 diode
R3303 N3302 N3303 10
D3303 N3303 0 diode
R3304 N3303 N3304 10
D3304 N3304 0 diode
R3305 N3304 N3305 10
D3305 N3305 0 diode
R3306 N3305 N3306 10
D3306 N3306 0 diode
R3307 N3306 N3307 10
D3307 N3307 0 diode
R3308 N3307 N3308 10
D3308 N3308 0 diode
R3309 N3308 N3309 10
D3309 N3309 0 diode
R3310 N3309 N3310 10
D3310 N3310 0 diode
R3311 N3310 N3311 10
D3311 N3311 0 diode
R3312 N3311 N3312 10
D3312 N3312 0 diode
R3313 N3312 N3313 10
D3313 N3313 0 diode
R3314 N3313 N3314 10
D3314 N3314 0 diode
R3315 N3314 N3315 10
D3315 N3315 0 diode
R3316 N3315 N3316 10
D3316 N3316 0 diode
R3317 N3316 N3317 10
D3317 N3317 0 diode
R3318 N3317 N3318 10
D3318 N3318 0 diode
R3319 N3318 N3319 10
D3319 N3319 0 diode
R3320 N3319 N3320 10
D3320 N3320 0 diode
R3321 N3320 N3321 10
D3321 N3321 0 diode
R3322 N3321 N3322 10
D3322 N3322 0 diode
R3323 N3322 N3323 10
D3323 N3323 0 diode
R3324 N3323 N3324 10
D3324 N3324 0 diode
R3325 N3324 N3325 10
D3325 N3325 0 diode
R3326 N3325 N3326 10
D3326 N3326 0 diode
R3327 N3326 N3327 10
D3327 N3327 0 diode
R3328 N3327 N3328 10
D3328 N3328 0 diode
R3329 N3328 N3329 10
D3329 N3329 0 diode
R3330 N3329 N3330 10
D3330 N3330 0 diode
R3331 N3330 N3331 10
D3331 N3331 0 diode
R3332 N3331 N3332 10
D3332 N3332 0 diode
R3333 N3332 N3333 10
D3333 N3333 0 diode
R3334 N3333 N3334 10
D3334 N3334 0 diode
R3335 N3334 N3335 10
D3335 N3335 0 diode
R3336 N3335 N3336 10
D3336 N3336 0 diode
R3337 N3336 N3337 10
D3337 N3337 0 diode
R3338 N3337 N3338 10
D3338 N3338 0 diode
R3339 N3338 N3339 10
D3339 N3339 0 diode
R3340 N3339 N3340 10
D3340 N3340 0 diode
R3341 N3340 N3341 10
D3341 N3341 0 diode
R3342 N3341 N3342 10
D3342 N3342 0 diode
R3343 N3342 N3343 10
D3343 N3343 0 diode
R3344 N3343 N3344 10
D3344 N3344 0 diode
R3345 N3344 N3345 10
D3345 N3345 0 diode
R3346 N3345 N3346 10
D3346 N3346 0 diode
R3347 N3346 N3347 10
D3347 N3347 0 diode
R3348 N3347 N3348 10
D3348 N3348 0 diode
R3349 N3348 N3349 10
D3349 N3349 0 diode
R3350 N3349 N3350 10
D3350 N3350 0 diode
R3351 N3350 N3351 10
D3351 N3351 0 diode
R3352 N3351 N3352 10
D3352 N3352 0 diode
R3353 N3352 N3353 10
D3353 N3353 0 diode
R3354 N3353 N3354 10
D3354 N3354 0 diode
R3355 N3354 N3355 10
D3355 N3355 0 diode
R3356 N3355 N3356 10
D3356 N3356 0 diode
R3357 N3356 N3357 10
D3357 N3357 0 diode
R3358 N3357 N3358 10
D3358 N3358 0 diode
R3359 N3358 N3359 10
D3359 N3359 0 diode
R3360 N3359 N3360 10
D3360 N3360 0 diode
R3361 N3360 N3361 10
D3361 N3361 0 diode
R3362 N3361 N3362 10
D3362 N3362 0 diode
R3363 N3362 N3363 10
D3363 N3363 0 diode
R3364 N3363 N3364 10
D3364 N3364 0 diode
R3365 N3364 N3365 10
D3365 N3365 0 diode
R3366 N3365 N3366 10
D3366 N3366 0 diode
R3367 N3366 N3367 10
D3367 N3367 0 diode
R3368 N3367 N3368 10
D3368 N3368 0 diode
R3369 N3368 N3369 10
D3369 N3369 0 diode
R3370 N3369 N3370 10
D3370 N3370 0 diode
R3371 N3370 N3371 10
D3371 N3371 0 diode
R3372 N3371 N3372 10
D3372 N3372 0 diode
R3373 N3372 N3373 10
D3373 N3373 0 diode
R3374 N3373 N3374 10
D3374 N3374 0 diode
R3375 N3374 N3375 10
D3375 N3375 0 diode
R3376 N3375 N3376 10
D3376 N3376 0 diode
R3377 N3376 N3377 10
D3377 N3377 0 diode
R3378 N3377 N3378 10
D3378 N3378 0 diode
R3379 N3378 N3379 10
D3379 N3379 0 diode
R3380 N3379 N3380 10
D3380 N3380 0 diode
R3381 N3380 N3381 10
D3381 N3381 0 diode
R3382 N3381 N3382 10
D3382 N3382 0 diode
R3383 N3382 N3383 10
D3383 N3383 0 diode
R3384 N3383 N3384 10
D3384 N3384 0 diode
R3385 N3384 N3385 10
D3385 N3385 0 diode
R3386 N3385 N3386 10
D3386 N3386 0 diode
R3387 N3386 N3387 10
D3387 N3387 0 diode
R3388 N3387 N3388 10
D3388 N3388 0 diode
R3389 N3388 N3389 10
D3389 N3389 0 diode
R3390 N3389 N3390 10
D3390 N3390 0 diode
R3391 N3390 N3391 10
D3391 N3391 0 diode
R3392 N3391 N3392 10
D3392 N3392 0 diode
R3393 N3392 N3393 10
D3393 N3393 0 diode
R3394 N3393 N3394 10
D3394 N3394 0 diode
R3395 N3394 N3395 10
D3395 N3395 0 diode
R3396 N3395 N3396 10
D3396 N3396 0 diode
R3397 N3396 N3397 10
D3397 N3397 0 diode
R3398 N3397 N3398 10
D3398 N3398 0 diode
R3399 N3398 N3399 10
D3399 N3399 0 diode
R3400 N3399 N3400 10
D3400 N3400 0 diode
R3401 N3400 N3401 10
D3401 N3401 0 diode
R3402 N3401 N3402 10
D3402 N3402 0 diode
R3403 N3402 N3403 10
D3403 N3403 0 diode
R3404 N3403 N3404 10
D3404 N3404 0 diode
R3405 N3404 N3405 10
D3405 N3405 0 diode
R3406 N3405 N3406 10
D3406 N3406 0 diode
R3407 N3406 N3407 10
D3407 N3407 0 diode
R3408 N3407 N3408 10
D3408 N3408 0 diode
R3409 N3408 N3409 10
D3409 N3409 0 diode
R3410 N3409 N3410 10
D3410 N3410 0 diode
R3411 N3410 N3411 10
D3411 N3411 0 diode
R3412 N3411 N3412 10
D3412 N3412 0 diode
R3413 N3412 N3413 10
D3413 N3413 0 diode
R3414 N3413 N3414 10
D3414 N3414 0 diode
R3415 N3414 N3415 10
D3415 N3415 0 diode
R3416 N3415 N3416 10
D3416 N3416 0 diode
R3417 N3416 N3417 10
D3417 N3417 0 diode
R3418 N3417 N3418 10
D3418 N3418 0 diode
R3419 N3418 N3419 10
D3419 N3419 0 diode
R3420 N3419 N3420 10
D3420 N3420 0 diode
R3421 N3420 N3421 10
D3421 N3421 0 diode
R3422 N3421 N3422 10
D3422 N3422 0 diode
R3423 N3422 N3423 10
D3423 N3423 0 diode
R3424 N3423 N3424 10
D3424 N3424 0 diode
R3425 N3424 N3425 10
D3425 N3425 0 diode
R3426 N3425 N3426 10
D3426 N3426 0 diode
R3427 N3426 N3427 10
D3427 N3427 0 diode
R3428 N3427 N3428 10
D3428 N3428 0 diode
R3429 N3428 N3429 10
D3429 N3429 0 diode
R3430 N3429 N3430 10
D3430 N3430 0 diode
R3431 N3430 N3431 10
D3431 N3431 0 diode
R3432 N3431 N3432 10
D3432 N3432 0 diode
R3433 N3432 N3433 10
D3433 N3433 0 diode
R3434 N3433 N3434 10
D3434 N3434 0 diode
R3435 N3434 N3435 10
D3435 N3435 0 diode
R3436 N3435 N3436 10
D3436 N3436 0 diode
R3437 N3436 N3437 10
D3437 N3437 0 diode
R3438 N3437 N3438 10
D3438 N3438 0 diode
R3439 N3438 N3439 10
D3439 N3439 0 diode
R3440 N3439 N3440 10
D3440 N3440 0 diode
R3441 N3440 N3441 10
D3441 N3441 0 diode
R3442 N3441 N3442 10
D3442 N3442 0 diode
R3443 N3442 N3443 10
D3443 N3443 0 diode
R3444 N3443 N3444 10
D3444 N3444 0 diode
R3445 N3444 N3445 10
D3445 N3445 0 diode
R3446 N3445 N3446 10
D3446 N3446 0 diode
R3447 N3446 N3447 10
D3447 N3447 0 diode
R3448 N3447 N3448 10
D3448 N3448 0 diode
R3449 N3448 N3449 10
D3449 N3449 0 diode
R3450 N3449 N3450 10
D3450 N3450 0 diode
R3451 N3450 N3451 10
D3451 N3451 0 diode
R3452 N3451 N3452 10
D3452 N3452 0 diode
R3453 N3452 N3453 10
D3453 N3453 0 diode
R3454 N3453 N3454 10
D3454 N3454 0 diode
R3455 N3454 N3455 10
D3455 N3455 0 diode
R3456 N3455 N3456 10
D3456 N3456 0 diode
R3457 N3456 N3457 10
D3457 N3457 0 diode
R3458 N3457 N3458 10
D3458 N3458 0 diode
R3459 N3458 N3459 10
D3459 N3459 0 diode
R3460 N3459 N3460 10
D3460 N3460 0 diode
R3461 N3460 N3461 10
D3461 N3461 0 diode
R3462 N3461 N3462 10
D3462 N3462 0 diode
R3463 N3462 N3463 10
D3463 N3463 0 diode
R3464 N3463 N3464 10
D3464 N3464 0 diode
R3465 N3464 N3465 10
D3465 N3465 0 diode
R3466 N3465 N3466 10
D3466 N3466 0 diode
R3467 N3466 N3467 10
D3467 N3467 0 diode
R3468 N3467 N3468 10
D3468 N3468 0 diode
R3469 N3468 N3469 10
D3469 N3469 0 diode
R3470 N3469 N3470 10
D3470 N3470 0 diode
R3471 N3470 N3471 10
D3471 N3471 0 diode
R3472 N3471 N3472 10
D3472 N3472 0 diode
R3473 N3472 N3473 10
D3473 N3473 0 diode
R3474 N3473 N3474 10
D3474 N3474 0 diode
R3475 N3474 N3475 10
D3475 N3475 0 diode
R3476 N3475 N3476 10
D3476 N3476 0 diode
R3477 N3476 N3477 10
D3477 N3477 0 diode
R3478 N3477 N3478 10
D3478 N3478 0 diode
R3479 N3478 N3479 10
D3479 N3479 0 diode
R3480 N3479 N3480 10
D3480 N3480 0 diode
R3481 N3480 N3481 10
D3481 N3481 0 diode
R3482 N3481 N3482 10
D3482 N3482 0 diode
R3483 N3482 N3483 10
D3483 N3483 0 diode
R3484 N3483 N3484 10
D3484 N3484 0 diode
R3485 N3484 N3485 10
D3485 N3485 0 diode
R3486 N3485 N3486 10
D3486 N3486 0 diode
R3487 N3486 N3487 10
D3487 N3487 0 diode
R3488 N3487 N3488 10
D3488 N3488 0 diode
R3489 N3488 N3489 10
D3489 N3489 0 diode
R3490 N3489 N3490 10
D3490 N3490 0 diode
R3491 N3490 N3491 10
D3491 N3491 0 diode
R3492 N3491 N3492 10
D3492 N3492 0 diode
R3493 N3492 N3493 10
D3493 N3493 0 diode
R3494 N3493 N3494 10
D3494 N3494 0 diode
R3495 N3494 N3495 10
D3495 N3495 0 diode
R3496 N3495 N3496 10
D3496 N3496 0 diode
R3497 N3496 N3497 10
D3497 N3497 0 diode
R3498 N3497 N3498 10
D3498 N3498 0 diode
R3499 N3498 N3499 10
D3499 N3499 0 diode
R3500 N3499 N3500 10
D3500 N3500 0 diode
R3501 N3500 N3501 10
D3501 N3501 0 diode
R3502 N3501 N3502 10
D3502 N3502 0 diode
R3503 N3502 N3503 10
D3503 N3503 0 diode
R3504 N3503 N3504 10
D3504 N3504 0 diode
R3505 N3504 N3505 10
D3505 N3505 0 diode
R3506 N3505 N3506 10
D3506 N3506 0 diode
R3507 N3506 N3507 10
D3507 N3507 0 diode
R3508 N3507 N3508 10
D3508 N3508 0 diode
R3509 N3508 N3509 10
D3509 N3509 0 diode
R3510 N3509 N3510 10
D3510 N3510 0 diode
R3511 N3510 N3511 10
D3511 N3511 0 diode
R3512 N3511 N3512 10
D3512 N3512 0 diode
R3513 N3512 N3513 10
D3513 N3513 0 diode
R3514 N3513 N3514 10
D3514 N3514 0 diode
R3515 N3514 N3515 10
D3515 N3515 0 diode
R3516 N3515 N3516 10
D3516 N3516 0 diode
R3517 N3516 N3517 10
D3517 N3517 0 diode
R3518 N3517 N3518 10
D3518 N3518 0 diode
R3519 N3518 N3519 10
D3519 N3519 0 diode
R3520 N3519 N3520 10
D3520 N3520 0 diode
R3521 N3520 N3521 10
D3521 N3521 0 diode
R3522 N3521 N3522 10
D3522 N3522 0 diode
R3523 N3522 N3523 10
D3523 N3523 0 diode
R3524 N3523 N3524 10
D3524 N3524 0 diode
R3525 N3524 N3525 10
D3525 N3525 0 diode
R3526 N3525 N3526 10
D3526 N3526 0 diode
R3527 N3526 N3527 10
D3527 N3527 0 diode
R3528 N3527 N3528 10
D3528 N3528 0 diode
R3529 N3528 N3529 10
D3529 N3529 0 diode
R3530 N3529 N3530 10
D3530 N3530 0 diode
R3531 N3530 N3531 10
D3531 N3531 0 diode
R3532 N3531 N3532 10
D3532 N3532 0 diode
R3533 N3532 N3533 10
D3533 N3533 0 diode
R3534 N3533 N3534 10
D3534 N3534 0 diode
R3535 N3534 N3535 10
D3535 N3535 0 diode
R3536 N3535 N3536 10
D3536 N3536 0 diode
R3537 N3536 N3537 10
D3537 N3537 0 diode
R3538 N3537 N3538 10
D3538 N3538 0 diode
R3539 N3538 N3539 10
D3539 N3539 0 diode
R3540 N3539 N3540 10
D3540 N3540 0 diode
R3541 N3540 N3541 10
D3541 N3541 0 diode
R3542 N3541 N3542 10
D3542 N3542 0 diode
R3543 N3542 N3543 10
D3543 N3543 0 diode
R3544 N3543 N3544 10
D3544 N3544 0 diode
R3545 N3544 N3545 10
D3545 N3545 0 diode
R3546 N3545 N3546 10
D3546 N3546 0 diode
R3547 N3546 N3547 10
D3547 N3547 0 diode
R3548 N3547 N3548 10
D3548 N3548 0 diode
R3549 N3548 N3549 10
D3549 N3549 0 diode
R3550 N3549 N3550 10
D3550 N3550 0 diode
R3551 N3550 N3551 10
D3551 N3551 0 diode
R3552 N3551 N3552 10
D3552 N3552 0 diode
R3553 N3552 N3553 10
D3553 N3553 0 diode
R3554 N3553 N3554 10
D3554 N3554 0 diode
R3555 N3554 N3555 10
D3555 N3555 0 diode
R3556 N3555 N3556 10
D3556 N3556 0 diode
R3557 N3556 N3557 10
D3557 N3557 0 diode
R3558 N3557 N3558 10
D3558 N3558 0 diode
R3559 N3558 N3559 10
D3559 N3559 0 diode
R3560 N3559 N3560 10
D3560 N3560 0 diode
R3561 N3560 N3561 10
D3561 N3561 0 diode
R3562 N3561 N3562 10
D3562 N3562 0 diode
R3563 N3562 N3563 10
D3563 N3563 0 diode
R3564 N3563 N3564 10
D3564 N3564 0 diode
R3565 N3564 N3565 10
D3565 N3565 0 diode
R3566 N3565 N3566 10
D3566 N3566 0 diode
R3567 N3566 N3567 10
D3567 N3567 0 diode
R3568 N3567 N3568 10
D3568 N3568 0 diode
R3569 N3568 N3569 10
D3569 N3569 0 diode
R3570 N3569 N3570 10
D3570 N3570 0 diode
R3571 N3570 N3571 10
D3571 N3571 0 diode
R3572 N3571 N3572 10
D3572 N3572 0 diode
R3573 N3572 N3573 10
D3573 N3573 0 diode
R3574 N3573 N3574 10
D3574 N3574 0 diode
R3575 N3574 N3575 10
D3575 N3575 0 diode
R3576 N3575 N3576 10
D3576 N3576 0 diode
R3577 N3576 N3577 10
D3577 N3577 0 diode
R3578 N3577 N3578 10
D3578 N3578 0 diode
R3579 N3578 N3579 10
D3579 N3579 0 diode
R3580 N3579 N3580 10
D3580 N3580 0 diode
R3581 N3580 N3581 10
D3581 N3581 0 diode
R3582 N3581 N3582 10
D3582 N3582 0 diode
R3583 N3582 N3583 10
D3583 N3583 0 diode
R3584 N3583 N3584 10
D3584 N3584 0 diode
R3585 N3584 N3585 10
D3585 N3585 0 diode
R3586 N3585 N3586 10
D3586 N3586 0 diode
R3587 N3586 N3587 10
D3587 N3587 0 diode
R3588 N3587 N3588 10
D3588 N3588 0 diode
R3589 N3588 N3589 10
D3589 N3589 0 diode
R3590 N3589 N3590 10
D3590 N3590 0 diode
R3591 N3590 N3591 10
D3591 N3591 0 diode
R3592 N3591 N3592 10
D3592 N3592 0 diode
R3593 N3592 N3593 10
D3593 N3593 0 diode
R3594 N3593 N3594 10
D3594 N3594 0 diode
R3595 N3594 N3595 10
D3595 N3595 0 diode
R3596 N3595 N3596 10
D3596 N3596 0 diode
R3597 N3596 N3597 10
D3597 N3597 0 diode
R3598 N3597 N3598 10
D3598 N3598 0 diode
R3599 N3598 N3599 10
D3599 N3599 0 diode
R3600 N3599 N3600 10
D3600 N3600 0 diode
R3601 N3600 N3601 10
D3601 N3601 0 diode
R3602 N3601 N3602 10
D3602 N3602 0 diode
R3603 N3602 N3603 10
D3603 N3603 0 diode
R3604 N3603 N3604 10
D3604 N3604 0 diode
R3605 N3604 N3605 10
D3605 N3605 0 diode
R3606 N3605 N3606 10
D3606 N3606 0 diode
R3607 N3606 N3607 10
D3607 N3607 0 diode
R3608 N3607 N3608 10
D3608 N3608 0 diode
R3609 N3608 N3609 10
D3609 N3609 0 diode
R3610 N3609 N3610 10
D3610 N3610 0 diode
R3611 N3610 N3611 10
D3611 N3611 0 diode
R3612 N3611 N3612 10
D3612 N3612 0 diode
R3613 N3612 N3613 10
D3613 N3613 0 diode
R3614 N3613 N3614 10
D3614 N3614 0 diode
R3615 N3614 N3615 10
D3615 N3615 0 diode
R3616 N3615 N3616 10
D3616 N3616 0 diode
R3617 N3616 N3617 10
D3617 N3617 0 diode
R3618 N3617 N3618 10
D3618 N3618 0 diode
R3619 N3618 N3619 10
D3619 N3619 0 diode
R3620 N3619 N3620 10
D3620 N3620 0 diode
R3621 N3620 N3621 10
D3621 N3621 0 diode
R3622 N3621 N3622 10
D3622 N3622 0 diode
R3623 N3622 N3623 10
D3623 N3623 0 diode
R3624 N3623 N3624 10
D3624 N3624 0 diode
R3625 N3624 N3625 10
D3625 N3625 0 diode
R3626 N3625 N3626 10
D3626 N3626 0 diode
R3627 N3626 N3627 10
D3627 N3627 0 diode
R3628 N3627 N3628 10
D3628 N3628 0 diode
R3629 N3628 N3629 10
D3629 N3629 0 diode
R3630 N3629 N3630 10
D3630 N3630 0 diode
R3631 N3630 N3631 10
D3631 N3631 0 diode
R3632 N3631 N3632 10
D3632 N3632 0 diode
R3633 N3632 N3633 10
D3633 N3633 0 diode
R3634 N3633 N3634 10
D3634 N3634 0 diode
R3635 N3634 N3635 10
D3635 N3635 0 diode
R3636 N3635 N3636 10
D3636 N3636 0 diode
R3637 N3636 N3637 10
D3637 N3637 0 diode
R3638 N3637 N3638 10
D3638 N3638 0 diode
R3639 N3638 N3639 10
D3639 N3639 0 diode
R3640 N3639 N3640 10
D3640 N3640 0 diode
R3641 N3640 N3641 10
D3641 N3641 0 diode
R3642 N3641 N3642 10
D3642 N3642 0 diode
R3643 N3642 N3643 10
D3643 N3643 0 diode
R3644 N3643 N3644 10
D3644 N3644 0 diode
R3645 N3644 N3645 10
D3645 N3645 0 diode
R3646 N3645 N3646 10
D3646 N3646 0 diode
R3647 N3646 N3647 10
D3647 N3647 0 diode
R3648 N3647 N3648 10
D3648 N3648 0 diode
R3649 N3648 N3649 10
D3649 N3649 0 diode
R3650 N3649 N3650 10
D3650 N3650 0 diode
R3651 N3650 N3651 10
D3651 N3651 0 diode
R3652 N3651 N3652 10
D3652 N3652 0 diode
R3653 N3652 N3653 10
D3653 N3653 0 diode
R3654 N3653 N3654 10
D3654 N3654 0 diode
R3655 N3654 N3655 10
D3655 N3655 0 diode
R3656 N3655 N3656 10
D3656 N3656 0 diode
R3657 N3656 N3657 10
D3657 N3657 0 diode
R3658 N3657 N3658 10
D3658 N3658 0 diode
R3659 N3658 N3659 10
D3659 N3659 0 diode
R3660 N3659 N3660 10
D3660 N3660 0 diode
R3661 N3660 N3661 10
D3661 N3661 0 diode
R3662 N3661 N3662 10
D3662 N3662 0 diode
R3663 N3662 N3663 10
D3663 N3663 0 diode
R3664 N3663 N3664 10
D3664 N3664 0 diode
R3665 N3664 N3665 10
D3665 N3665 0 diode
R3666 N3665 N3666 10
D3666 N3666 0 diode
R3667 N3666 N3667 10
D3667 N3667 0 diode
R3668 N3667 N3668 10
D3668 N3668 0 diode
R3669 N3668 N3669 10
D3669 N3669 0 diode
R3670 N3669 N3670 10
D3670 N3670 0 diode
R3671 N3670 N3671 10
D3671 N3671 0 diode
R3672 N3671 N3672 10
D3672 N3672 0 diode
R3673 N3672 N3673 10
D3673 N3673 0 diode
R3674 N3673 N3674 10
D3674 N3674 0 diode
R3675 N3674 N3675 10
D3675 N3675 0 diode
R3676 N3675 N3676 10
D3676 N3676 0 diode
R3677 N3676 N3677 10
D3677 N3677 0 diode
R3678 N3677 N3678 10
D3678 N3678 0 diode
R3679 N3678 N3679 10
D3679 N3679 0 diode
R3680 N3679 N3680 10
D3680 N3680 0 diode
R3681 N3680 N3681 10
D3681 N3681 0 diode
R3682 N3681 N3682 10
D3682 N3682 0 diode
R3683 N3682 N3683 10
D3683 N3683 0 diode
R3684 N3683 N3684 10
D3684 N3684 0 diode
R3685 N3684 N3685 10
D3685 N3685 0 diode
R3686 N3685 N3686 10
D3686 N3686 0 diode
R3687 N3686 N3687 10
D3687 N3687 0 diode
R3688 N3687 N3688 10
D3688 N3688 0 diode
R3689 N3688 N3689 10
D3689 N3689 0 diode
R3690 N3689 N3690 10
D3690 N3690 0 diode
R3691 N3690 N3691 10
D3691 N3691 0 diode
R3692 N3691 N3692 10
D3692 N3692 0 diode
R3693 N3692 N3693 10
D3693 N3693 0 diode
R3694 N3693 N3694 10
D3694 N3694 0 diode
R3695 N3694 N3695 10
D3695 N3695 0 diode
R3696 N3695 N3696 10
D3696 N3696 0 diode
R3697 N3696 N3697 10
D3697 N3697 0 diode
R3698 N3697 N3698 10
D3698 N3698 0 diode
R3699 N3698 N3699 10
D3699 N3699 0 diode
R3700 N3699 N3700 10
D3700 N3700 0 diode
R3701 N3700 N3701 10
D3701 N3701 0 diode
R3702 N3701 N3702 10
D3702 N3702 0 diode
R3703 N3702 N3703 10
D3703 N3703 0 diode
R3704 N3703 N3704 10
D3704 N3704 0 diode
R3705 N3704 N3705 10
D3705 N3705 0 diode
R3706 N3705 N3706 10
D3706 N3706 0 diode
R3707 N3706 N3707 10
D3707 N3707 0 diode
R3708 N3707 N3708 10
D3708 N3708 0 diode
R3709 N3708 N3709 10
D3709 N3709 0 diode
R3710 N3709 N3710 10
D3710 N3710 0 diode
R3711 N3710 N3711 10
D3711 N3711 0 diode
R3712 N3711 N3712 10
D3712 N3712 0 diode
R3713 N3712 N3713 10
D3713 N3713 0 diode
R3714 N3713 N3714 10
D3714 N3714 0 diode
R3715 N3714 N3715 10
D3715 N3715 0 diode
R3716 N3715 N3716 10
D3716 N3716 0 diode
R3717 N3716 N3717 10
D3717 N3717 0 diode
R3718 N3717 N3718 10
D3718 N3718 0 diode
R3719 N3718 N3719 10
D3719 N3719 0 diode
R3720 N3719 N3720 10
D3720 N3720 0 diode
R3721 N3720 N3721 10
D3721 N3721 0 diode
R3722 N3721 N3722 10
D3722 N3722 0 diode
R3723 N3722 N3723 10
D3723 N3723 0 diode
R3724 N3723 N3724 10
D3724 N3724 0 diode
R3725 N3724 N3725 10
D3725 N3725 0 diode
R3726 N3725 N3726 10
D3726 N3726 0 diode
R3727 N3726 N3727 10
D3727 N3727 0 diode
R3728 N3727 N3728 10
D3728 N3728 0 diode
R3729 N3728 N3729 10
D3729 N3729 0 diode
R3730 N3729 N3730 10
D3730 N3730 0 diode
R3731 N3730 N3731 10
D3731 N3731 0 diode
R3732 N3731 N3732 10
D3732 N3732 0 diode
R3733 N3732 N3733 10
D3733 N3733 0 diode
R3734 N3733 N3734 10
D3734 N3734 0 diode
R3735 N3734 N3735 10
D3735 N3735 0 diode
R3736 N3735 N3736 10
D3736 N3736 0 diode
R3737 N3736 N3737 10
D3737 N3737 0 diode
R3738 N3737 N3738 10
D3738 N3738 0 diode
R3739 N3738 N3739 10
D3739 N3739 0 diode
R3740 N3739 N3740 10
D3740 N3740 0 diode
R3741 N3740 N3741 10
D3741 N3741 0 diode
R3742 N3741 N3742 10
D3742 N3742 0 diode
R3743 N3742 N3743 10
D3743 N3743 0 diode
R3744 N3743 N3744 10
D3744 N3744 0 diode
R3745 N3744 N3745 10
D3745 N3745 0 diode
R3746 N3745 N3746 10
D3746 N3746 0 diode
R3747 N3746 N3747 10
D3747 N3747 0 diode
R3748 N3747 N3748 10
D3748 N3748 0 diode
R3749 N3748 N3749 10
D3749 N3749 0 diode
R3750 N3749 N3750 10
D3750 N3750 0 diode
R3751 N3750 N3751 10
D3751 N3751 0 diode
R3752 N3751 N3752 10
D3752 N3752 0 diode
R3753 N3752 N3753 10
D3753 N3753 0 diode
R3754 N3753 N3754 10
D3754 N3754 0 diode
R3755 N3754 N3755 10
D3755 N3755 0 diode
R3756 N3755 N3756 10
D3756 N3756 0 diode
R3757 N3756 N3757 10
D3757 N3757 0 diode
R3758 N3757 N3758 10
D3758 N3758 0 diode
R3759 N3758 N3759 10
D3759 N3759 0 diode
R3760 N3759 N3760 10
D3760 N3760 0 diode
R3761 N3760 N3761 10
D3761 N3761 0 diode
R3762 N3761 N3762 10
D3762 N3762 0 diode
R3763 N3762 N3763 10
D3763 N3763 0 diode
R3764 N3763 N3764 10
D3764 N3764 0 diode
R3765 N3764 N3765 10
D3765 N3765 0 diode
R3766 N3765 N3766 10
D3766 N3766 0 diode
R3767 N3766 N3767 10
D3767 N3767 0 diode
R3768 N3767 N3768 10
D3768 N3768 0 diode
R3769 N3768 N3769 10
D3769 N3769 0 diode
R3770 N3769 N3770 10
D3770 N3770 0 diode
R3771 N3770 N3771 10
D3771 N3771 0 diode
R3772 N3771 N3772 10
D3772 N3772 0 diode
R3773 N3772 N3773 10
D3773 N3773 0 diode
R3774 N3773 N3774 10
D3774 N3774 0 diode
R3775 N3774 N3775 10
D3775 N3775 0 diode
R3776 N3775 N3776 10
D3776 N3776 0 diode
R3777 N3776 N3777 10
D3777 N3777 0 diode
R3778 N3777 N3778 10
D3778 N3778 0 diode
R3779 N3778 N3779 10
D3779 N3779 0 diode
R3780 N3779 N3780 10
D3780 N3780 0 diode
R3781 N3780 N3781 10
D3781 N3781 0 diode
R3782 N3781 N3782 10
D3782 N3782 0 diode
R3783 N3782 N3783 10
D3783 N3783 0 diode
R3784 N3783 N3784 10
D3784 N3784 0 diode
R3785 N3784 N3785 10
D3785 N3785 0 diode
R3786 N3785 N3786 10
D3786 N3786 0 diode
R3787 N3786 N3787 10
D3787 N3787 0 diode
R3788 N3787 N3788 10
D3788 N3788 0 diode
R3789 N3788 N3789 10
D3789 N3789 0 diode
R3790 N3789 N3790 10
D3790 N3790 0 diode
R3791 N3790 N3791 10
D3791 N3791 0 diode
R3792 N3791 N3792 10
D3792 N3792 0 diode
R3793 N3792 N3793 10
D3793 N3793 0 diode
R3794 N3793 N3794 10
D3794 N3794 0 diode
R3795 N3794 N3795 10
D3795 N3795 0 diode
R3796 N3795 N3796 10
D3796 N3796 0 diode
R3797 N3796 N3797 10
D3797 N3797 0 diode
R3798 N3797 N3798 10
D3798 N3798 0 diode
R3799 N3798 N3799 10
D3799 N3799 0 diode
R3800 N3799 N3800 10
D3800 N3800 0 diode
R3801 N3800 N3801 10
D3801 N3801 0 diode
R3802 N3801 N3802 10
D3802 N3802 0 diode
R3803 N3802 N3803 10
D3803 N3803 0 diode
R3804 N3803 N3804 10
D3804 N3804 0 diode
R3805 N3804 N3805 10
D3805 N3805 0 diode
R3806 N3805 N3806 10
D3806 N3806 0 diode
R3807 N3806 N3807 10
D3807 N3807 0 diode
R3808 N3807 N3808 10
D3808 N3808 0 diode
R3809 N3808 N3809 10
D3809 N3809 0 diode
R3810 N3809 N3810 10
D3810 N3810 0 diode
R3811 N3810 N3811 10
D3811 N3811 0 diode
R3812 N3811 N3812 10
D3812 N3812 0 diode
R3813 N3812 N3813 10
D3813 N3813 0 diode
R3814 N3813 N3814 10
D3814 N3814 0 diode
R3815 N3814 N3815 10
D3815 N3815 0 diode
R3816 N3815 N3816 10
D3816 N3816 0 diode
R3817 N3816 N3817 10
D3817 N3817 0 diode
R3818 N3817 N3818 10
D3818 N3818 0 diode
R3819 N3818 N3819 10
D3819 N3819 0 diode
R3820 N3819 N3820 10
D3820 N3820 0 diode
R3821 N3820 N3821 10
D3821 N3821 0 diode
R3822 N3821 N3822 10
D3822 N3822 0 diode
R3823 N3822 N3823 10
D3823 N3823 0 diode
R3824 N3823 N3824 10
D3824 N3824 0 diode
R3825 N3824 N3825 10
D3825 N3825 0 diode
R3826 N3825 N3826 10
D3826 N3826 0 diode
R3827 N3826 N3827 10
D3827 N3827 0 diode
R3828 N3827 N3828 10
D3828 N3828 0 diode
R3829 N3828 N3829 10
D3829 N3829 0 diode
R3830 N3829 N3830 10
D3830 N3830 0 diode
R3831 N3830 N3831 10
D3831 N3831 0 diode
R3832 N3831 N3832 10
D3832 N3832 0 diode
R3833 N3832 N3833 10
D3833 N3833 0 diode
R3834 N3833 N3834 10
D3834 N3834 0 diode
R3835 N3834 N3835 10
D3835 N3835 0 diode
R3836 N3835 N3836 10
D3836 N3836 0 diode
R3837 N3836 N3837 10
D3837 N3837 0 diode
R3838 N3837 N3838 10
D3838 N3838 0 diode
R3839 N3838 N3839 10
D3839 N3839 0 diode
R3840 N3839 N3840 10
D3840 N3840 0 diode
R3841 N3840 N3841 10
D3841 N3841 0 diode
R3842 N3841 N3842 10
D3842 N3842 0 diode
R3843 N3842 N3843 10
D3843 N3843 0 diode
R3844 N3843 N3844 10
D3844 N3844 0 diode
R3845 N3844 N3845 10
D3845 N3845 0 diode
R3846 N3845 N3846 10
D3846 N3846 0 diode
R3847 N3846 N3847 10
D3847 N3847 0 diode
R3848 N3847 N3848 10
D3848 N3848 0 diode
R3849 N3848 N3849 10
D3849 N3849 0 diode
R3850 N3849 N3850 10
D3850 N3850 0 diode
R3851 N3850 N3851 10
D3851 N3851 0 diode
R3852 N3851 N3852 10
D3852 N3852 0 diode
R3853 N3852 N3853 10
D3853 N3853 0 diode
R3854 N3853 N3854 10
D3854 N3854 0 diode
R3855 N3854 N3855 10
D3855 N3855 0 diode
R3856 N3855 N3856 10
D3856 N3856 0 diode
R3857 N3856 N3857 10
D3857 N3857 0 diode
R3858 N3857 N3858 10
D3858 N3858 0 diode
R3859 N3858 N3859 10
D3859 N3859 0 diode
R3860 N3859 N3860 10
D3860 N3860 0 diode
R3861 N3860 N3861 10
D3861 N3861 0 diode
R3862 N3861 N3862 10
D3862 N3862 0 diode
R3863 N3862 N3863 10
D3863 N3863 0 diode
R3864 N3863 N3864 10
D3864 N3864 0 diode
R3865 N3864 N3865 10
D3865 N3865 0 diode
R3866 N3865 N3866 10
D3866 N3866 0 diode
R3867 N3866 N3867 10
D3867 N3867 0 diode
R3868 N3867 N3868 10
D3868 N3868 0 diode
R3869 N3868 N3869 10
D3869 N3869 0 diode
R3870 N3869 N3870 10
D3870 N3870 0 diode
R3871 N3870 N3871 10
D3871 N3871 0 diode
R3872 N3871 N3872 10
D3872 N3872 0 diode
R3873 N3872 N3873 10
D3873 N3873 0 diode
R3874 N3873 N3874 10
D3874 N3874 0 diode
R3875 N3874 N3875 10
D3875 N3875 0 diode
R3876 N3875 N3876 10
D3876 N3876 0 diode
R3877 N3876 N3877 10
D3877 N3877 0 diode
R3878 N3877 N3878 10
D3878 N3878 0 diode
R3879 N3878 N3879 10
D3879 N3879 0 diode
R3880 N3879 N3880 10
D3880 N3880 0 diode
R3881 N3880 N3881 10
D3881 N3881 0 diode
R3882 N3881 N3882 10
D3882 N3882 0 diode
R3883 N3882 N3883 10
D3883 N3883 0 diode
R3884 N3883 N3884 10
D3884 N3884 0 diode
R3885 N3884 N3885 10
D3885 N3885 0 diode
R3886 N3885 N3886 10
D3886 N3886 0 diode
R3887 N3886 N3887 10
D3887 N3887 0 diode
R3888 N3887 N3888 10
D3888 N3888 0 diode
R3889 N3888 N3889 10
D3889 N3889 0 diode
R3890 N3889 N3890 10
D3890 N3890 0 diode
R3891 N3890 N3891 10
D3891 N3891 0 diode
R3892 N3891 N3892 10
D3892 N3892 0 diode
R3893 N3892 N3893 10
D3893 N3893 0 diode
R3894 N3893 N3894 10
D3894 N3894 0 diode
R3895 N3894 N3895 10
D3895 N3895 0 diode
R3896 N3895 N3896 10
D3896 N3896 0 diode
R3897 N3896 N3897 10
D3897 N3897 0 diode
R3898 N3897 N3898 10
D3898 N3898 0 diode
R3899 N3898 N3899 10
D3899 N3899 0 diode
R3900 N3899 N3900 10
D3900 N3900 0 diode
R3901 N3900 N3901 10
D3901 N3901 0 diode
R3902 N3901 N3902 10
D3902 N3902 0 diode
R3903 N3902 N3903 10
D3903 N3903 0 diode
R3904 N3903 N3904 10
D3904 N3904 0 diode
R3905 N3904 N3905 10
D3905 N3905 0 diode
R3906 N3905 N3906 10
D3906 N3906 0 diode
R3907 N3906 N3907 10
D3907 N3907 0 diode
R3908 N3907 N3908 10
D3908 N3908 0 diode
R3909 N3908 N3909 10
D3909 N3909 0 diode
R3910 N3909 N3910 10
D3910 N3910 0 diode
R3911 N3910 N3911 10
D3911 N3911 0 diode
R3912 N3911 N3912 10
D3912 N3912 0 diode
R3913 N3912 N3913 10
D3913 N3913 0 diode
R3914 N3913 N3914 10
D3914 N3914 0 diode
R3915 N3914 N3915 10
D3915 N3915 0 diode
R3916 N3915 N3916 10
D3916 N3916 0 diode
R3917 N3916 N3917 10
D3917 N3917 0 diode
R3918 N3917 N3918 10
D3918 N3918 0 diode
R3919 N3918 N3919 10
D3919 N3919 0 diode
R3920 N3919 N3920 10
D3920 N3920 0 diode
R3921 N3920 N3921 10
D3921 N3921 0 diode
R3922 N3921 N3922 10
D3922 N3922 0 diode
R3923 N3922 N3923 10
D3923 N3923 0 diode
R3924 N3923 N3924 10
D3924 N3924 0 diode
R3925 N3924 N3925 10
D3925 N3925 0 diode
R3926 N3925 N3926 10
D3926 N3926 0 diode
R3927 N3926 N3927 10
D3927 N3927 0 diode
R3928 N3927 N3928 10
D3928 N3928 0 diode
R3929 N3928 N3929 10
D3929 N3929 0 diode
R3930 N3929 N3930 10
D3930 N3930 0 diode
R3931 N3930 N3931 10
D3931 N3931 0 diode
R3932 N3931 N3932 10
D3932 N3932 0 diode
R3933 N3932 N3933 10
D3933 N3933 0 diode
R3934 N3933 N3934 10
D3934 N3934 0 diode
R3935 N3934 N3935 10
D3935 N3935 0 diode
R3936 N3935 N3936 10
D3936 N3936 0 diode
R3937 N3936 N3937 10
D3937 N3937 0 diode
R3938 N3937 N3938 10
D3938 N3938 0 diode
R3939 N3938 N3939 10
D3939 N3939 0 diode
R3940 N3939 N3940 10
D3940 N3940 0 diode
R3941 N3940 N3941 10
D3941 N3941 0 diode
R3942 N3941 N3942 10
D3942 N3942 0 diode
R3943 N3942 N3943 10
D3943 N3943 0 diode
R3944 N3943 N3944 10
D3944 N3944 0 diode
R3945 N3944 N3945 10
D3945 N3945 0 diode
R3946 N3945 N3946 10
D3946 N3946 0 diode
R3947 N3946 N3947 10
D3947 N3947 0 diode
R3948 N3947 N3948 10
D3948 N3948 0 diode
R3949 N3948 N3949 10
D3949 N3949 0 diode
R3950 N3949 N3950 10
D3950 N3950 0 diode
R3951 N3950 N3951 10
D3951 N3951 0 diode
R3952 N3951 N3952 10
D3952 N3952 0 diode
R3953 N3952 N3953 10
D3953 N3953 0 diode
R3954 N3953 N3954 10
D3954 N3954 0 diode
R3955 N3954 N3955 10
D3955 N3955 0 diode
R3956 N3955 N3956 10
D3956 N3956 0 diode
R3957 N3956 N3957 10
D3957 N3957 0 diode
R3958 N3957 N3958 10
D3958 N3958 0 diode
R3959 N3958 N3959 10
D3959 N3959 0 diode
R3960 N3959 N3960 10
D3960 N3960 0 diode
R3961 N3960 N3961 10
D3961 N3961 0 diode
R3962 N3961 N3962 10
D3962 N3962 0 diode
R3963 N3962 N3963 10
D3963 N3963 0 diode
R3964 N3963 N3964 10
D3964 N3964 0 diode
R3965 N3964 N3965 10
D3965 N3965 0 diode
R3966 N3965 N3966 10
D3966 N3966 0 diode
R3967 N3966 N3967 10
D3967 N3967 0 diode
R3968 N3967 N3968 10
D3968 N3968 0 diode
R3969 N3968 N3969 10
D3969 N3969 0 diode
R3970 N3969 N3970 10
D3970 N3970 0 diode
R3971 N3970 N3971 10
D3971 N3971 0 diode
R3972 N3971 N3972 10
D3972 N3972 0 diode
R3973 N3972 N3973 10
D3973 N3973 0 diode
R3974 N3973 N3974 10
D3974 N3974 0 diode
R3975 N3974 N3975 10
D3975 N3975 0 diode
R3976 N3975 N3976 10
D3976 N3976 0 diode
R3977 N3976 N3977 10
D3977 N3977 0 diode
R3978 N3977 N3978 10
D3978 N3978 0 diode
R3979 N3978 N3979 10
D3979 N3979 0 diode
R3980 N3979 N3980 10
D3980 N3980 0 diode
R3981 N3980 N3981 10
D3981 N3981 0 diode
R3982 N3981 N3982 10
D3982 N3982 0 diode
R3983 N3982 N3983 10
D3983 N3983 0 diode
R3984 N3983 N3984 10
D3984 N3984 0 diode
R3985 N3984 N3985 10
D3985 N3985 0 diode
R3986 N3985 N3986 10
D3986 N3986 0 diode
R3987 N3986 N3987 10
D3987 N3987 0 diode
R3988 N3987 N3988 10
D3988 N3988 0 diode
R3989 N3988 N3989 10
D3989 N3989 0 diode
R3990 N3989 N3990 10
D3990 N3990 0 diode
R3991 N3990 N3991 10
D3991 N3991 0 diode
R3992 N3991 N3992 10
D3992 N3992 0 diode
R3993 N3992 N3993 10
D3993 N3993 0 diode
R3994 N3993 N3994 10
D3994 N3994 0 diode
R3995 N3994 N3995 10
D3995 N3995 0 diode
R3996 N3995 N3996 10
D3996 N3996 0 diode
R3997 N3996 N3997 10
D3997 N3997 0 diode
R3998 N3997 N3998 10
D3998 N3998 0 diode
R3999 N3998 N3999 10
D3999 N3999 0 diode
R4000 N3999 N4000 10
D4000 N4000 0 diode
R4001 N4000 N4001 10
D4001 N4001 0 diode
R4002 N4001 N4002 10
D4002 N4002 0 diode
R4003 N4002 N4003 10
D4003 N4003 0 diode
R4004 N4003 N4004 10
D4004 N4004 0 diode
R4005 N4004 N4005 10
D4005 N4005 0 diode
R4006 N4005 N4006 10
D4006 N4006 0 diode
R4007 N4006 N4007 10
D4007 N4007 0 diode
R4008 N4007 N4008 10
D4008 N4008 0 diode
R4009 N4008 N4009 10
D4009 N4009 0 diode
R4010 N4009 N4010 10
D4010 N4010 0 diode
R4011 N4010 N4011 10
D4011 N4011 0 diode
R4012 N4011 N4012 10
D4012 N4012 0 diode
R4013 N4012 N4013 10
D4013 N4013 0 diode
R4014 N4013 N4014 10
D4014 N4014 0 diode
R4015 N4014 N4015 10
D4015 N4015 0 diode
R4016 N4015 N4016 10
D4016 N4016 0 diode
R4017 N4016 N4017 10
D4017 N4017 0 diode
R4018 N4017 N4018 10
D4018 N4018 0 diode
R4019 N4018 N4019 10
D4019 N4019 0 diode
R4020 N4019 N4020 10
D4020 N4020 0 diode
R4021 N4020 N4021 10
D4021 N4021 0 diode
R4022 N4021 N4022 10
D4022 N4022 0 diode
R4023 N4022 N4023 10
D4023 N4023 0 diode
R4024 N4023 N4024 10
D4024 N4024 0 diode
R4025 N4024 N4025 10
D4025 N4025 0 diode
R4026 N4025 N4026 10
D4026 N4026 0 diode
R4027 N4026 N4027 10
D4027 N4027 0 diode
R4028 N4027 N4028 10
D4028 N4028 0 diode
R4029 N4028 N4029 10
D4029 N4029 0 diode
R4030 N4029 N4030 10
D4030 N4030 0 diode
R4031 N4030 N4031 10
D4031 N4031 0 diode
R4032 N4031 N4032 10
D4032 N4032 0 diode
R4033 N4032 N4033 10
D4033 N4033 0 diode
R4034 N4033 N4034 10
D4034 N4034 0 diode
R4035 N4034 N4035 10
D4035 N4035 0 diode
R4036 N4035 N4036 10
D4036 N4036 0 diode
R4037 N4036 N4037 10
D4037 N4037 0 diode
R4038 N4037 N4038 10
D4038 N4038 0 diode
R4039 N4038 N4039 10
D4039 N4039 0 diode
R4040 N4039 N4040 10
D4040 N4040 0 diode
R4041 N4040 N4041 10
D4041 N4041 0 diode
R4042 N4041 N4042 10
D4042 N4042 0 diode
R4043 N4042 N4043 10
D4043 N4043 0 diode
R4044 N4043 N4044 10
D4044 N4044 0 diode
R4045 N4044 N4045 10
D4045 N4045 0 diode
R4046 N4045 N4046 10
D4046 N4046 0 diode
R4047 N4046 N4047 10
D4047 N4047 0 diode
R4048 N4047 N4048 10
D4048 N4048 0 diode
R4049 N4048 N4049 10
D4049 N4049 0 diode
R4050 N4049 N4050 10
D4050 N4050 0 diode
R4051 N4050 N4051 10
D4051 N4051 0 diode
R4052 N4051 N4052 10
D4052 N4052 0 diode
R4053 N4052 N4053 10
D4053 N4053 0 diode
R4054 N4053 N4054 10
D4054 N4054 0 diode
R4055 N4054 N4055 10
D4055 N4055 0 diode
R4056 N4055 N4056 10
D4056 N4056 0 diode
R4057 N4056 N4057 10
D4057 N4057 0 diode
R4058 N4057 N4058 10
D4058 N4058 0 diode
R4059 N4058 N4059 10
D4059 N4059 0 diode
R4060 N4059 N4060 10
D4060 N4060 0 diode
R4061 N4060 N4061 10
D4061 N4061 0 diode
R4062 N4061 N4062 10
D4062 N4062 0 diode
R4063 N4062 N4063 10
D4063 N4063 0 diode
R4064 N4063 N4064 10
D4064 N4064 0 diode
R4065 N4064 N4065 10
D4065 N4065 0 diode
R4066 N4065 N4066 10
D4066 N4066 0 diode
R4067 N4066 N4067 10
D4067 N4067 0 diode
R4068 N4067 N4068 10
D4068 N4068 0 diode
R4069 N4068 N4069 10
D4069 N4069 0 diode
R4070 N4069 N4070 10
D4070 N4070 0 diode
R4071 N4070 N4071 10
D4071 N4071 0 diode
R4072 N4071 N4072 10
D4072 N4072 0 diode
R4073 N4072 N4073 10
D4073 N4073 0 diode
R4074 N4073 N4074 10
D4074 N4074 0 diode
R4075 N4074 N4075 10
D4075 N4075 0 diode
R4076 N4075 N4076 10
D4076 N4076 0 diode
R4077 N4076 N4077 10
D4077 N4077 0 diode
R4078 N4077 N4078 10
D4078 N4078 0 diode
R4079 N4078 N4079 10
D4079 N4079 0 diode
R4080 N4079 N4080 10
D4080 N4080 0 diode
R4081 N4080 N4081 10
D4081 N4081 0 diode
R4082 N4081 N4082 10
D4082 N4082 0 diode
R4083 N4082 N4083 10
D4083 N4083 0 diode
R4084 N4083 N4084 10
D4084 N4084 0 diode
R4085 N4084 N4085 10
D4085 N4085 0 diode
R4086 N4085 N4086 10
D4086 N4086 0 diode
R4087 N4086 N4087 10
D4087 N4087 0 diode
R4088 N4087 N4088 10
D4088 N4088 0 diode
R4089 N4088 N4089 10
D4089 N4089 0 diode
R4090 N4089 N4090 10
D4090 N4090 0 diode
R4091 N4090 N4091 10
D4091 N4091 0 diode
R4092 N4091 N4092 10
D4092 N4092 0 diode
R4093 N4092 N4093 10
D4093 N4093 0 diode
R4094 N4093 N4094 10
D4094 N4094 0 diode
R4095 N4094 N4095 10
D4095 N4095 0 diode
R4096 N4095 N4096 10
D4096 N4096 0 diode
R4097 N4096 N4097 10
D4097 N4097 0 diode
R4098 N4097 N4098 10
D4098 N4098 0 diode
R4099 N4098 N4099 10
D4099 N4099 0 diode
R4100 N4099 N4100 10
D4100 N4100 0 diode
R4101 N4100 N4101 10
D4101 N4101 0 diode
R4102 N4101 N4102 10
D4102 N4102 0 diode
R4103 N4102 N4103 10
D4103 N4103 0 diode
R4104 N4103 N4104 10
D4104 N4104 0 diode
R4105 N4104 N4105 10
D4105 N4105 0 diode
R4106 N4105 N4106 10
D4106 N4106 0 diode
R4107 N4106 N4107 10
D4107 N4107 0 diode
R4108 N4107 N4108 10
D4108 N4108 0 diode
R4109 N4108 N4109 10
D4109 N4109 0 diode
R4110 N4109 N4110 10
D4110 N4110 0 diode
R4111 N4110 N4111 10
D4111 N4111 0 diode
R4112 N4111 N4112 10
D4112 N4112 0 diode
R4113 N4112 N4113 10
D4113 N4113 0 diode
R4114 N4113 N4114 10
D4114 N4114 0 diode
R4115 N4114 N4115 10
D4115 N4115 0 diode
R4116 N4115 N4116 10
D4116 N4116 0 diode
R4117 N4116 N4117 10
D4117 N4117 0 diode
R4118 N4117 N4118 10
D4118 N4118 0 diode
R4119 N4118 N4119 10
D4119 N4119 0 diode
R4120 N4119 N4120 10
D4120 N4120 0 diode
R4121 N4120 N4121 10
D4121 N4121 0 diode
R4122 N4121 N4122 10
D4122 N4122 0 diode
R4123 N4122 N4123 10
D4123 N4123 0 diode
R4124 N4123 N4124 10
D4124 N4124 0 diode
R4125 N4124 N4125 10
D4125 N4125 0 diode
R4126 N4125 N4126 10
D4126 N4126 0 diode
R4127 N4126 N4127 10
D4127 N4127 0 diode
R4128 N4127 N4128 10
D4128 N4128 0 diode
R4129 N4128 N4129 10
D4129 N4129 0 diode
R4130 N4129 N4130 10
D4130 N4130 0 diode
R4131 N4130 N4131 10
D4131 N4131 0 diode
R4132 N4131 N4132 10
D4132 N4132 0 diode
R4133 N4132 N4133 10
D4133 N4133 0 diode
R4134 N4133 N4134 10
D4134 N4134 0 diode
R4135 N4134 N4135 10
D4135 N4135 0 diode
R4136 N4135 N4136 10
D4136 N4136 0 diode
R4137 N4136 N4137 10
D4137 N4137 0 diode
R4138 N4137 N4138 10
D4138 N4138 0 diode
R4139 N4138 N4139 10
D4139 N4139 0 diode
R4140 N4139 N4140 10
D4140 N4140 0 diode
R4141 N4140 N4141 10
D4141 N4141 0 diode
R4142 N4141 N4142 10
D4142 N4142 0 diode
R4143 N4142 N4143 10
D4143 N4143 0 diode
R4144 N4143 N4144 10
D4144 N4144 0 diode
R4145 N4144 N4145 10
D4145 N4145 0 diode
R4146 N4145 N4146 10
D4146 N4146 0 diode
R4147 N4146 N4147 10
D4147 N4147 0 diode
R4148 N4147 N4148 10
D4148 N4148 0 diode
R4149 N4148 N4149 10
D4149 N4149 0 diode
R4150 N4149 N4150 10
D4150 N4150 0 diode
R4151 N4150 N4151 10
D4151 N4151 0 diode
R4152 N4151 N4152 10
D4152 N4152 0 diode
R4153 N4152 N4153 10
D4153 N4153 0 diode
R4154 N4153 N4154 10
D4154 N4154 0 diode
R4155 N4154 N4155 10
D4155 N4155 0 diode
R4156 N4155 N4156 10
D4156 N4156 0 diode
R4157 N4156 N4157 10
D4157 N4157 0 diode
R4158 N4157 N4158 10
D4158 N4158 0 diode
R4159 N4158 N4159 10
D4159 N4159 0 diode
R4160 N4159 N4160 10
D4160 N4160 0 diode
R4161 N4160 N4161 10
D4161 N4161 0 diode
R4162 N4161 N4162 10
D4162 N4162 0 diode
R4163 N4162 N4163 10
D4163 N4163 0 diode
R4164 N4163 N4164 10
D4164 N4164 0 diode
R4165 N4164 N4165 10
D4165 N4165 0 diode
R4166 N4165 N4166 10
D4166 N4166 0 diode
R4167 N4166 N4167 10
D4167 N4167 0 diode
R4168 N4167 N4168 10
D4168 N4168 0 diode
R4169 N4168 N4169 10
D4169 N4169 0 diode
R4170 N4169 N4170 10
D4170 N4170 0 diode
R4171 N4170 N4171 10
D4171 N4171 0 diode
R4172 N4171 N4172 10
D4172 N4172 0 diode
R4173 N4172 N4173 10
D4173 N4173 0 diode
R4174 N4173 N4174 10
D4174 N4174 0 diode
R4175 N4174 N4175 10
D4175 N4175 0 diode
R4176 N4175 N4176 10
D4176 N4176 0 diode
R4177 N4176 N4177 10
D4177 N4177 0 diode
R4178 N4177 N4178 10
D4178 N4178 0 diode
R4179 N4178 N4179 10
D4179 N4179 0 diode
R4180 N4179 N4180 10
D4180 N4180 0 diode
R4181 N4180 N4181 10
D4181 N4181 0 diode
R4182 N4181 N4182 10
D4182 N4182 0 diode
R4183 N4182 N4183 10
D4183 N4183 0 diode
R4184 N4183 N4184 10
D4184 N4184 0 diode
R4185 N4184 N4185 10
D4185 N4185 0 diode
R4186 N4185 N4186 10
D4186 N4186 0 diode
R4187 N4186 N4187 10
D4187 N4187 0 diode
R4188 N4187 N4188 10
D4188 N4188 0 diode
R4189 N4188 N4189 10
D4189 N4189 0 diode
R4190 N4189 N4190 10
D4190 N4190 0 diode
R4191 N4190 N4191 10
D4191 N4191 0 diode
R4192 N4191 N4192 10
D4192 N4192 0 diode
R4193 N4192 N4193 10
D4193 N4193 0 diode
R4194 N4193 N4194 10
D4194 N4194 0 diode
R4195 N4194 N4195 10
D4195 N4195 0 diode
R4196 N4195 N4196 10
D4196 N4196 0 diode
R4197 N4196 N4197 10
D4197 N4197 0 diode
R4198 N4197 N4198 10
D4198 N4198 0 diode
R4199 N4198 N4199 10
D4199 N4199 0 diode
R4200 N4199 N4200 10
D4200 N4200 0 diode
R4201 N4200 N4201 10
D4201 N4201 0 diode
R4202 N4201 N4202 10
D4202 N4202 0 diode
R4203 N4202 N4203 10
D4203 N4203 0 diode
R4204 N4203 N4204 10
D4204 N4204 0 diode
R4205 N4204 N4205 10
D4205 N4205 0 diode
R4206 N4205 N4206 10
D4206 N4206 0 diode
R4207 N4206 N4207 10
D4207 N4207 0 diode
R4208 N4207 N4208 10
D4208 N4208 0 diode
R4209 N4208 N4209 10
D4209 N4209 0 diode
R4210 N4209 N4210 10
D4210 N4210 0 diode
R4211 N4210 N4211 10
D4211 N4211 0 diode
R4212 N4211 N4212 10
D4212 N4212 0 diode
R4213 N4212 N4213 10
D4213 N4213 0 diode
R4214 N4213 N4214 10
D4214 N4214 0 diode
R4215 N4214 N4215 10
D4215 N4215 0 diode
R4216 N4215 N4216 10
D4216 N4216 0 diode
R4217 N4216 N4217 10
D4217 N4217 0 diode
R4218 N4217 N4218 10
D4218 N4218 0 diode
R4219 N4218 N4219 10
D4219 N4219 0 diode
R4220 N4219 N4220 10
D4220 N4220 0 diode
R4221 N4220 N4221 10
D4221 N4221 0 diode
R4222 N4221 N4222 10
D4222 N4222 0 diode
R4223 N4222 N4223 10
D4223 N4223 0 diode
R4224 N4223 N4224 10
D4224 N4224 0 diode
R4225 N4224 N4225 10
D4225 N4225 0 diode
R4226 N4225 N4226 10
D4226 N4226 0 diode
R4227 N4226 N4227 10
D4227 N4227 0 diode
R4228 N4227 N4228 10
D4228 N4228 0 diode
R4229 N4228 N4229 10
D4229 N4229 0 diode
R4230 N4229 N4230 10
D4230 N4230 0 diode
R4231 N4230 N4231 10
D4231 N4231 0 diode
R4232 N4231 N4232 10
D4232 N4232 0 diode
R4233 N4232 N4233 10
D4233 N4233 0 diode
R4234 N4233 N4234 10
D4234 N4234 0 diode
R4235 N4234 N4235 10
D4235 N4235 0 diode
R4236 N4235 N4236 10
D4236 N4236 0 diode
R4237 N4236 N4237 10
D4237 N4237 0 diode
R4238 N4237 N4238 10
D4238 N4238 0 diode
R4239 N4238 N4239 10
D4239 N4239 0 diode
R4240 N4239 N4240 10
D4240 N4240 0 diode
R4241 N4240 N4241 10
D4241 N4241 0 diode
R4242 N4241 N4242 10
D4242 N4242 0 diode
R4243 N4242 N4243 10
D4243 N4243 0 diode
R4244 N4243 N4244 10
D4244 N4244 0 diode
R4245 N4244 N4245 10
D4245 N4245 0 diode
R4246 N4245 N4246 10
D4246 N4246 0 diode
R4247 N4246 N4247 10
D4247 N4247 0 diode
R4248 N4247 N4248 10
D4248 N4248 0 diode
R4249 N4248 N4249 10
D4249 N4249 0 diode
R4250 N4249 N4250 10
D4250 N4250 0 diode
R4251 N4250 N4251 10
D4251 N4251 0 diode
R4252 N4251 N4252 10
D4252 N4252 0 diode
R4253 N4252 N4253 10
D4253 N4253 0 diode
R4254 N4253 N4254 10
D4254 N4254 0 diode
R4255 N4254 N4255 10
D4255 N4255 0 diode
R4256 N4255 N4256 10
D4256 N4256 0 diode
R4257 N4256 N4257 10
D4257 N4257 0 diode
R4258 N4257 N4258 10
D4258 N4258 0 diode
R4259 N4258 N4259 10
D4259 N4259 0 diode
R4260 N4259 N4260 10
D4260 N4260 0 diode
R4261 N4260 N4261 10
D4261 N4261 0 diode
R4262 N4261 N4262 10
D4262 N4262 0 diode
R4263 N4262 N4263 10
D4263 N4263 0 diode
R4264 N4263 N4264 10
D4264 N4264 0 diode
R4265 N4264 N4265 10
D4265 N4265 0 diode
R4266 N4265 N4266 10
D4266 N4266 0 diode
R4267 N4266 N4267 10
D4267 N4267 0 diode
R4268 N4267 N4268 10
D4268 N4268 0 diode
R4269 N4268 N4269 10
D4269 N4269 0 diode
R4270 N4269 N4270 10
D4270 N4270 0 diode
R4271 N4270 N4271 10
D4271 N4271 0 diode
R4272 N4271 N4272 10
D4272 N4272 0 diode
R4273 N4272 N4273 10
D4273 N4273 0 diode
R4274 N4273 N4274 10
D4274 N4274 0 diode
R4275 N4274 N4275 10
D4275 N4275 0 diode
R4276 N4275 N4276 10
D4276 N4276 0 diode
R4277 N4276 N4277 10
D4277 N4277 0 diode
R4278 N4277 N4278 10
D4278 N4278 0 diode
R4279 N4278 N4279 10
D4279 N4279 0 diode
R4280 N4279 N4280 10
D4280 N4280 0 diode
R4281 N4280 N4281 10
D4281 N4281 0 diode
R4282 N4281 N4282 10
D4282 N4282 0 diode
R4283 N4282 N4283 10
D4283 N4283 0 diode
R4284 N4283 N4284 10
D4284 N4284 0 diode
R4285 N4284 N4285 10
D4285 N4285 0 diode
R4286 N4285 N4286 10
D4286 N4286 0 diode
R4287 N4286 N4287 10
D4287 N4287 0 diode
R4288 N4287 N4288 10
D4288 N4288 0 diode
R4289 N4288 N4289 10
D4289 N4289 0 diode
R4290 N4289 N4290 10
D4290 N4290 0 diode
R4291 N4290 N4291 10
D4291 N4291 0 diode
R4292 N4291 N4292 10
D4292 N4292 0 diode
R4293 N4292 N4293 10
D4293 N4293 0 diode
R4294 N4293 N4294 10
D4294 N4294 0 diode
R4295 N4294 N4295 10
D4295 N4295 0 diode
R4296 N4295 N4296 10
D4296 N4296 0 diode
R4297 N4296 N4297 10
D4297 N4297 0 diode
R4298 N4297 N4298 10
D4298 N4298 0 diode
R4299 N4298 N4299 10
D4299 N4299 0 diode
R4300 N4299 N4300 10
D4300 N4300 0 diode
R4301 N4300 N4301 10
D4301 N4301 0 diode
R4302 N4301 N4302 10
D4302 N4302 0 diode
R4303 N4302 N4303 10
D4303 N4303 0 diode
R4304 N4303 N4304 10
D4304 N4304 0 diode
R4305 N4304 N4305 10
D4305 N4305 0 diode
R4306 N4305 N4306 10
D4306 N4306 0 diode
R4307 N4306 N4307 10
D4307 N4307 0 diode
R4308 N4307 N4308 10
D4308 N4308 0 diode
R4309 N4308 N4309 10
D4309 N4309 0 diode
R4310 N4309 N4310 10
D4310 N4310 0 diode
R4311 N4310 N4311 10
D4311 N4311 0 diode
R4312 N4311 N4312 10
D4312 N4312 0 diode
R4313 N4312 N4313 10
D4313 N4313 0 diode
R4314 N4313 N4314 10
D4314 N4314 0 diode
R4315 N4314 N4315 10
D4315 N4315 0 diode
R4316 N4315 N4316 10
D4316 N4316 0 diode
R4317 N4316 N4317 10
D4317 N4317 0 diode
R4318 N4317 N4318 10
D4318 N4318 0 diode
R4319 N4318 N4319 10
D4319 N4319 0 diode
R4320 N4319 N4320 10
D4320 N4320 0 diode
R4321 N4320 N4321 10
D4321 N4321 0 diode
R4322 N4321 N4322 10
D4322 N4322 0 diode
R4323 N4322 N4323 10
D4323 N4323 0 diode
R4324 N4323 N4324 10
D4324 N4324 0 diode
R4325 N4324 N4325 10
D4325 N4325 0 diode
R4326 N4325 N4326 10
D4326 N4326 0 diode
R4327 N4326 N4327 10
D4327 N4327 0 diode
R4328 N4327 N4328 10
D4328 N4328 0 diode
R4329 N4328 N4329 10
D4329 N4329 0 diode
R4330 N4329 N4330 10
D4330 N4330 0 diode
R4331 N4330 N4331 10
D4331 N4331 0 diode
R4332 N4331 N4332 10
D4332 N4332 0 diode
R4333 N4332 N4333 10
D4333 N4333 0 diode
R4334 N4333 N4334 10
D4334 N4334 0 diode
R4335 N4334 N4335 10
D4335 N4335 0 diode
R4336 N4335 N4336 10
D4336 N4336 0 diode
R4337 N4336 N4337 10
D4337 N4337 0 diode
R4338 N4337 N4338 10
D4338 N4338 0 diode
R4339 N4338 N4339 10
D4339 N4339 0 diode
R4340 N4339 N4340 10
D4340 N4340 0 diode
R4341 N4340 N4341 10
D4341 N4341 0 diode
R4342 N4341 N4342 10
D4342 N4342 0 diode
R4343 N4342 N4343 10
D4343 N4343 0 diode
R4344 N4343 N4344 10
D4344 N4344 0 diode
R4345 N4344 N4345 10
D4345 N4345 0 diode
R4346 N4345 N4346 10
D4346 N4346 0 diode
R4347 N4346 N4347 10
D4347 N4347 0 diode
R4348 N4347 N4348 10
D4348 N4348 0 diode
R4349 N4348 N4349 10
D4349 N4349 0 diode
R4350 N4349 N4350 10
D4350 N4350 0 diode
R4351 N4350 N4351 10
D4351 N4351 0 diode
R4352 N4351 N4352 10
D4352 N4352 0 diode
R4353 N4352 N4353 10
D4353 N4353 0 diode
R4354 N4353 N4354 10
D4354 N4354 0 diode
R4355 N4354 N4355 10
D4355 N4355 0 diode
R4356 N4355 N4356 10
D4356 N4356 0 diode
R4357 N4356 N4357 10
D4357 N4357 0 diode
R4358 N4357 N4358 10
D4358 N4358 0 diode
R4359 N4358 N4359 10
D4359 N4359 0 diode
R4360 N4359 N4360 10
D4360 N4360 0 diode
R4361 N4360 N4361 10
D4361 N4361 0 diode
R4362 N4361 N4362 10
D4362 N4362 0 diode
R4363 N4362 N4363 10
D4363 N4363 0 diode
R4364 N4363 N4364 10
D4364 N4364 0 diode
R4365 N4364 N4365 10
D4365 N4365 0 diode
R4366 N4365 N4366 10
D4366 N4366 0 diode
R4367 N4366 N4367 10
D4367 N4367 0 diode
R4368 N4367 N4368 10
D4368 N4368 0 diode
R4369 N4368 N4369 10
D4369 N4369 0 diode
R4370 N4369 N4370 10
D4370 N4370 0 diode
R4371 N4370 N4371 10
D4371 N4371 0 diode
R4372 N4371 N4372 10
D4372 N4372 0 diode
R4373 N4372 N4373 10
D4373 N4373 0 diode
R4374 N4373 N4374 10
D4374 N4374 0 diode
R4375 N4374 N4375 10
D4375 N4375 0 diode
R4376 N4375 N4376 10
D4376 N4376 0 diode
R4377 N4376 N4377 10
D4377 N4377 0 diode
R4378 N4377 N4378 10
D4378 N4378 0 diode
R4379 N4378 N4379 10
D4379 N4379 0 diode
R4380 N4379 N4380 10
D4380 N4380 0 diode
R4381 N4380 N4381 10
D4381 N4381 0 diode
R4382 N4381 N4382 10
D4382 N4382 0 diode
R4383 N4382 N4383 10
D4383 N4383 0 diode
R4384 N4383 N4384 10
D4384 N4384 0 diode
R4385 N4384 N4385 10
D4385 N4385 0 diode
R4386 N4385 N4386 10
D4386 N4386 0 diode
R4387 N4386 N4387 10
D4387 N4387 0 diode
R4388 N4387 N4388 10
D4388 N4388 0 diode
R4389 N4388 N4389 10
D4389 N4389 0 diode
R4390 N4389 N4390 10
D4390 N4390 0 diode
R4391 N4390 N4391 10
D4391 N4391 0 diode
R4392 N4391 N4392 10
D4392 N4392 0 diode
R4393 N4392 N4393 10
D4393 N4393 0 diode
R4394 N4393 N4394 10
D4394 N4394 0 diode
R4395 N4394 N4395 10
D4395 N4395 0 diode
R4396 N4395 N4396 10
D4396 N4396 0 diode
R4397 N4396 N4397 10
D4397 N4397 0 diode
R4398 N4397 N4398 10
D4398 N4398 0 diode
R4399 N4398 N4399 10
D4399 N4399 0 diode
R4400 N4399 N4400 10
D4400 N4400 0 diode
R4401 N4400 N4401 10
D4401 N4401 0 diode
R4402 N4401 N4402 10
D4402 N4402 0 diode
R4403 N4402 N4403 10
D4403 N4403 0 diode
R4404 N4403 N4404 10
D4404 N4404 0 diode
R4405 N4404 N4405 10
D4405 N4405 0 diode
R4406 N4405 N4406 10
D4406 N4406 0 diode
R4407 N4406 N4407 10
D4407 N4407 0 diode
R4408 N4407 N4408 10
D4408 N4408 0 diode
R4409 N4408 N4409 10
D4409 N4409 0 diode
R4410 N4409 N4410 10
D4410 N4410 0 diode
R4411 N4410 N4411 10
D4411 N4411 0 diode
R4412 N4411 N4412 10
D4412 N4412 0 diode
R4413 N4412 N4413 10
D4413 N4413 0 diode
R4414 N4413 N4414 10
D4414 N4414 0 diode
R4415 N4414 N4415 10
D4415 N4415 0 diode
R4416 N4415 N4416 10
D4416 N4416 0 diode
R4417 N4416 N4417 10
D4417 N4417 0 diode
R4418 N4417 N4418 10
D4418 N4418 0 diode
R4419 N4418 N4419 10
D4419 N4419 0 diode
R4420 N4419 N4420 10
D4420 N4420 0 diode
R4421 N4420 N4421 10
D4421 N4421 0 diode
R4422 N4421 N4422 10
D4422 N4422 0 diode
R4423 N4422 N4423 10
D4423 N4423 0 diode
R4424 N4423 N4424 10
D4424 N4424 0 diode
R4425 N4424 N4425 10
D4425 N4425 0 diode
R4426 N4425 N4426 10
D4426 N4426 0 diode
R4427 N4426 N4427 10
D4427 N4427 0 diode
R4428 N4427 N4428 10
D4428 N4428 0 diode
R4429 N4428 N4429 10
D4429 N4429 0 diode
R4430 N4429 N4430 10
D4430 N4430 0 diode
R4431 N4430 N4431 10
D4431 N4431 0 diode
R4432 N4431 N4432 10
D4432 N4432 0 diode
R4433 N4432 N4433 10
D4433 N4433 0 diode
R4434 N4433 N4434 10
D4434 N4434 0 diode
R4435 N4434 N4435 10
D4435 N4435 0 diode
R4436 N4435 N4436 10
D4436 N4436 0 diode
R4437 N4436 N4437 10
D4437 N4437 0 diode
R4438 N4437 N4438 10
D4438 N4438 0 diode
R4439 N4438 N4439 10
D4439 N4439 0 diode
R4440 N4439 N4440 10
D4440 N4440 0 diode
R4441 N4440 N4441 10
D4441 N4441 0 diode
R4442 N4441 N4442 10
D4442 N4442 0 diode
R4443 N4442 N4443 10
D4443 N4443 0 diode
R4444 N4443 N4444 10
D4444 N4444 0 diode
R4445 N4444 N4445 10
D4445 N4445 0 diode
R4446 N4445 N4446 10
D4446 N4446 0 diode
R4447 N4446 N4447 10
D4447 N4447 0 diode
R4448 N4447 N4448 10
D4448 N4448 0 diode
R4449 N4448 N4449 10
D4449 N4449 0 diode
R4450 N4449 N4450 10
D4450 N4450 0 diode
R4451 N4450 N4451 10
D4451 N4451 0 diode
R4452 N4451 N4452 10
D4452 N4452 0 diode
R4453 N4452 N4453 10
D4453 N4453 0 diode
R4454 N4453 N4454 10
D4454 N4454 0 diode
R4455 N4454 N4455 10
D4455 N4455 0 diode
R4456 N4455 N4456 10
D4456 N4456 0 diode
R4457 N4456 N4457 10
D4457 N4457 0 diode
R4458 N4457 N4458 10
D4458 N4458 0 diode
R4459 N4458 N4459 10
D4459 N4459 0 diode
R4460 N4459 N4460 10
D4460 N4460 0 diode
R4461 N4460 N4461 10
D4461 N4461 0 diode
R4462 N4461 N4462 10
D4462 N4462 0 diode
R4463 N4462 N4463 10
D4463 N4463 0 diode
R4464 N4463 N4464 10
D4464 N4464 0 diode
R4465 N4464 N4465 10
D4465 N4465 0 diode
R4466 N4465 N4466 10
D4466 N4466 0 diode
R4467 N4466 N4467 10
D4467 N4467 0 diode
R4468 N4467 N4468 10
D4468 N4468 0 diode
R4469 N4468 N4469 10
D4469 N4469 0 diode
R4470 N4469 N4470 10
D4470 N4470 0 diode
R4471 N4470 N4471 10
D4471 N4471 0 diode
R4472 N4471 N4472 10
D4472 N4472 0 diode
R4473 N4472 N4473 10
D4473 N4473 0 diode
R4474 N4473 N4474 10
D4474 N4474 0 diode
R4475 N4474 N4475 10
D4475 N4475 0 diode
R4476 N4475 N4476 10
D4476 N4476 0 diode
R4477 N4476 N4477 10
D4477 N4477 0 diode
R4478 N4477 N4478 10
D4478 N4478 0 diode
R4479 N4478 N4479 10
D4479 N4479 0 diode
R4480 N4479 N4480 10
D4480 N4480 0 diode
R4481 N4480 N4481 10
D4481 N4481 0 diode
R4482 N4481 N4482 10
D4482 N4482 0 diode
R4483 N4482 N4483 10
D4483 N4483 0 diode
R4484 N4483 N4484 10
D4484 N4484 0 diode
R4485 N4484 N4485 10
D4485 N4485 0 diode
R4486 N4485 N4486 10
D4486 N4486 0 diode
R4487 N4486 N4487 10
D4487 N4487 0 diode
R4488 N4487 N4488 10
D4488 N4488 0 diode
R4489 N4488 N4489 10
D4489 N4489 0 diode
R4490 N4489 N4490 10
D4490 N4490 0 diode
R4491 N4490 N4491 10
D4491 N4491 0 diode
R4492 N4491 N4492 10
D4492 N4492 0 diode
R4493 N4492 N4493 10
D4493 N4493 0 diode
R4494 N4493 N4494 10
D4494 N4494 0 diode
R4495 N4494 N4495 10
D4495 N4495 0 diode
R4496 N4495 N4496 10
D4496 N4496 0 diode
R4497 N4496 N4497 10
D4497 N4497 0 diode
R4498 N4497 N4498 10
D4498 N4498 0 diode
R4499 N4498 N4499 10
D4499 N4499 0 diode
R4500 N4499 N4500 10
D4500 N4500 0 diode
R4501 N4500 N4501 10
D4501 N4501 0 diode
R4502 N4501 N4502 10
D4502 N4502 0 diode
R4503 N4502 N4503 10
D4503 N4503 0 diode
R4504 N4503 N4504 10
D4504 N4504 0 diode
R4505 N4504 N4505 10
D4505 N4505 0 diode
R4506 N4505 N4506 10
D4506 N4506 0 diode
R4507 N4506 N4507 10
D4507 N4507 0 diode
R4508 N4507 N4508 10
D4508 N4508 0 diode
R4509 N4508 N4509 10
D4509 N4509 0 diode
R4510 N4509 N4510 10
D4510 N4510 0 diode
R4511 N4510 N4511 10
D4511 N4511 0 diode
R4512 N4511 N4512 10
D4512 N4512 0 diode
R4513 N4512 N4513 10
D4513 N4513 0 diode
R4514 N4513 N4514 10
D4514 N4514 0 diode
R4515 N4514 N4515 10
D4515 N4515 0 diode
R4516 N4515 N4516 10
D4516 N4516 0 diode
R4517 N4516 N4517 10
D4517 N4517 0 diode
R4518 N4517 N4518 10
D4518 N4518 0 diode
R4519 N4518 N4519 10
D4519 N4519 0 diode
R4520 N4519 N4520 10
D4520 N4520 0 diode
R4521 N4520 N4521 10
D4521 N4521 0 diode
R4522 N4521 N4522 10
D4522 N4522 0 diode
R4523 N4522 N4523 10
D4523 N4523 0 diode
R4524 N4523 N4524 10
D4524 N4524 0 diode
R4525 N4524 N4525 10
D4525 N4525 0 diode
R4526 N4525 N4526 10
D4526 N4526 0 diode
R4527 N4526 N4527 10
D4527 N4527 0 diode
R4528 N4527 N4528 10
D4528 N4528 0 diode
R4529 N4528 N4529 10
D4529 N4529 0 diode
R4530 N4529 N4530 10
D4530 N4530 0 diode
R4531 N4530 N4531 10
D4531 N4531 0 diode
R4532 N4531 N4532 10
D4532 N4532 0 diode
R4533 N4532 N4533 10
D4533 N4533 0 diode
R4534 N4533 N4534 10
D4534 N4534 0 diode
R4535 N4534 N4535 10
D4535 N4535 0 diode
R4536 N4535 N4536 10
D4536 N4536 0 diode
R4537 N4536 N4537 10
D4537 N4537 0 diode
R4538 N4537 N4538 10
D4538 N4538 0 diode
R4539 N4538 N4539 10
D4539 N4539 0 diode
R4540 N4539 N4540 10
D4540 N4540 0 diode
R4541 N4540 N4541 10
D4541 N4541 0 diode
R4542 N4541 N4542 10
D4542 N4542 0 diode
R4543 N4542 N4543 10
D4543 N4543 0 diode
R4544 N4543 N4544 10
D4544 N4544 0 diode
R4545 N4544 N4545 10
D4545 N4545 0 diode
R4546 N4545 N4546 10
D4546 N4546 0 diode
R4547 N4546 N4547 10
D4547 N4547 0 diode
R4548 N4547 N4548 10
D4548 N4548 0 diode
R4549 N4548 N4549 10
D4549 N4549 0 diode
R4550 N4549 N4550 10
D4550 N4550 0 diode
R4551 N4550 N4551 10
D4551 N4551 0 diode
R4552 N4551 N4552 10
D4552 N4552 0 diode
R4553 N4552 N4553 10
D4553 N4553 0 diode
R4554 N4553 N4554 10
D4554 N4554 0 diode
R4555 N4554 N4555 10
D4555 N4555 0 diode
R4556 N4555 N4556 10
D4556 N4556 0 diode
R4557 N4556 N4557 10
D4557 N4557 0 diode
R4558 N4557 N4558 10
D4558 N4558 0 diode
R4559 N4558 N4559 10
D4559 N4559 0 diode
R4560 N4559 N4560 10
D4560 N4560 0 diode
R4561 N4560 N4561 10
D4561 N4561 0 diode
R4562 N4561 N4562 10
D4562 N4562 0 diode
R4563 N4562 N4563 10
D4563 N4563 0 diode
R4564 N4563 N4564 10
D4564 N4564 0 diode
R4565 N4564 N4565 10
D4565 N4565 0 diode
R4566 N4565 N4566 10
D4566 N4566 0 diode
R4567 N4566 N4567 10
D4567 N4567 0 diode
R4568 N4567 N4568 10
D4568 N4568 0 diode
R4569 N4568 N4569 10
D4569 N4569 0 diode
R4570 N4569 N4570 10
D4570 N4570 0 diode
R4571 N4570 N4571 10
D4571 N4571 0 diode
R4572 N4571 N4572 10
D4572 N4572 0 diode
R4573 N4572 N4573 10
D4573 N4573 0 diode
R4574 N4573 N4574 10
D4574 N4574 0 diode
R4575 N4574 N4575 10
D4575 N4575 0 diode
R4576 N4575 N4576 10
D4576 N4576 0 diode
R4577 N4576 N4577 10
D4577 N4577 0 diode
R4578 N4577 N4578 10
D4578 N4578 0 diode
R4579 N4578 N4579 10
D4579 N4579 0 diode
R4580 N4579 N4580 10
D4580 N4580 0 diode
R4581 N4580 N4581 10
D4581 N4581 0 diode
R4582 N4581 N4582 10
D4582 N4582 0 diode
R4583 N4582 N4583 10
D4583 N4583 0 diode
R4584 N4583 N4584 10
D4584 N4584 0 diode
R4585 N4584 N4585 10
D4585 N4585 0 diode
R4586 N4585 N4586 10
D4586 N4586 0 diode
R4587 N4586 N4587 10
D4587 N4587 0 diode
R4588 N4587 N4588 10
D4588 N4588 0 diode
R4589 N4588 N4589 10
D4589 N4589 0 diode
R4590 N4589 N4590 10
D4590 N4590 0 diode
R4591 N4590 N4591 10
D4591 N4591 0 diode
R4592 N4591 N4592 10
D4592 N4592 0 diode
R4593 N4592 N4593 10
D4593 N4593 0 diode
R4594 N4593 N4594 10
D4594 N4594 0 diode
R4595 N4594 N4595 10
D4595 N4595 0 diode
R4596 N4595 N4596 10
D4596 N4596 0 diode
R4597 N4596 N4597 10
D4597 N4597 0 diode
R4598 N4597 N4598 10
D4598 N4598 0 diode
R4599 N4598 N4599 10
D4599 N4599 0 diode
R4600 N4599 N4600 10
D4600 N4600 0 diode
R4601 N4600 N4601 10
D4601 N4601 0 diode
R4602 N4601 N4602 10
D4602 N4602 0 diode
R4603 N4602 N4603 10
D4603 N4603 0 diode
R4604 N4603 N4604 10
D4604 N4604 0 diode
R4605 N4604 N4605 10
D4605 N4605 0 diode
R4606 N4605 N4606 10
D4606 N4606 0 diode
R4607 N4606 N4607 10
D4607 N4607 0 diode
R4608 N4607 N4608 10
D4608 N4608 0 diode
R4609 N4608 N4609 10
D4609 N4609 0 diode
R4610 N4609 N4610 10
D4610 N4610 0 diode
R4611 N4610 N4611 10
D4611 N4611 0 diode
R4612 N4611 N4612 10
D4612 N4612 0 diode
R4613 N4612 N4613 10
D4613 N4613 0 diode
R4614 N4613 N4614 10
D4614 N4614 0 diode
R4615 N4614 N4615 10
D4615 N4615 0 diode
R4616 N4615 N4616 10
D4616 N4616 0 diode
R4617 N4616 N4617 10
D4617 N4617 0 diode
R4618 N4617 N4618 10
D4618 N4618 0 diode
R4619 N4618 N4619 10
D4619 N4619 0 diode
R4620 N4619 N4620 10
D4620 N4620 0 diode
R4621 N4620 N4621 10
D4621 N4621 0 diode
R4622 N4621 N4622 10
D4622 N4622 0 diode
R4623 N4622 N4623 10
D4623 N4623 0 diode
R4624 N4623 N4624 10
D4624 N4624 0 diode
R4625 N4624 N4625 10
D4625 N4625 0 diode
R4626 N4625 N4626 10
D4626 N4626 0 diode
R4627 N4626 N4627 10
D4627 N4627 0 diode
R4628 N4627 N4628 10
D4628 N4628 0 diode
R4629 N4628 N4629 10
D4629 N4629 0 diode
R4630 N4629 N4630 10
D4630 N4630 0 diode
R4631 N4630 N4631 10
D4631 N4631 0 diode
R4632 N4631 N4632 10
D4632 N4632 0 diode
R4633 N4632 N4633 10
D4633 N4633 0 diode
R4634 N4633 N4634 10
D4634 N4634 0 diode
R4635 N4634 N4635 10
D4635 N4635 0 diode
R4636 N4635 N4636 10
D4636 N4636 0 diode
R4637 N4636 N4637 10
D4637 N4637 0 diode
R4638 N4637 N4638 10
D4638 N4638 0 diode
R4639 N4638 N4639 10
D4639 N4639 0 diode
R4640 N4639 N4640 10
D4640 N4640 0 diode
R4641 N4640 N4641 10
D4641 N4641 0 diode
R4642 N4641 N4642 10
D4642 N4642 0 diode
R4643 N4642 N4643 10
D4643 N4643 0 diode
R4644 N4643 N4644 10
D4644 N4644 0 diode
R4645 N4644 N4645 10
D4645 N4645 0 diode
R4646 N4645 N4646 10
D4646 N4646 0 diode
R4647 N4646 N4647 10
D4647 N4647 0 diode
R4648 N4647 N4648 10
D4648 N4648 0 diode
R4649 N4648 N4649 10
D4649 N4649 0 diode
R4650 N4649 N4650 10
D4650 N4650 0 diode
R4651 N4650 N4651 10
D4651 N4651 0 diode
R4652 N4651 N4652 10
D4652 N4652 0 diode
R4653 N4652 N4653 10
D4653 N4653 0 diode
R4654 N4653 N4654 10
D4654 N4654 0 diode
R4655 N4654 N4655 10
D4655 N4655 0 diode
R4656 N4655 N4656 10
D4656 N4656 0 diode
R4657 N4656 N4657 10
D4657 N4657 0 diode
R4658 N4657 N4658 10
D4658 N4658 0 diode
R4659 N4658 N4659 10
D4659 N4659 0 diode
R4660 N4659 N4660 10
D4660 N4660 0 diode
R4661 N4660 N4661 10
D4661 N4661 0 diode
R4662 N4661 N4662 10
D4662 N4662 0 diode
R4663 N4662 N4663 10
D4663 N4663 0 diode
R4664 N4663 N4664 10
D4664 N4664 0 diode
R4665 N4664 N4665 10
D4665 N4665 0 diode
R4666 N4665 N4666 10
D4666 N4666 0 diode
R4667 N4666 N4667 10
D4667 N4667 0 diode
R4668 N4667 N4668 10
D4668 N4668 0 diode
R4669 N4668 N4669 10
D4669 N4669 0 diode
R4670 N4669 N4670 10
D4670 N4670 0 diode
R4671 N4670 N4671 10
D4671 N4671 0 diode
R4672 N4671 N4672 10
D4672 N4672 0 diode
R4673 N4672 N4673 10
D4673 N4673 0 diode
R4674 N4673 N4674 10
D4674 N4674 0 diode
R4675 N4674 N4675 10
D4675 N4675 0 diode
R4676 N4675 N4676 10
D4676 N4676 0 diode
R4677 N4676 N4677 10
D4677 N4677 0 diode
R4678 N4677 N4678 10
D4678 N4678 0 diode
R4679 N4678 N4679 10
D4679 N4679 0 diode
R4680 N4679 N4680 10
D4680 N4680 0 diode
R4681 N4680 N4681 10
D4681 N4681 0 diode
R4682 N4681 N4682 10
D4682 N4682 0 diode
R4683 N4682 N4683 10
D4683 N4683 0 diode
R4684 N4683 N4684 10
D4684 N4684 0 diode
R4685 N4684 N4685 10
D4685 N4685 0 diode
R4686 N4685 N4686 10
D4686 N4686 0 diode
R4687 N4686 N4687 10
D4687 N4687 0 diode
R4688 N4687 N4688 10
D4688 N4688 0 diode
R4689 N4688 N4689 10
D4689 N4689 0 diode
R4690 N4689 N4690 10
D4690 N4690 0 diode
R4691 N4690 N4691 10
D4691 N4691 0 diode
R4692 N4691 N4692 10
D4692 N4692 0 diode
R4693 N4692 N4693 10
D4693 N4693 0 diode
R4694 N4693 N4694 10
D4694 N4694 0 diode
R4695 N4694 N4695 10
D4695 N4695 0 diode
R4696 N4695 N4696 10
D4696 N4696 0 diode
R4697 N4696 N4697 10
D4697 N4697 0 diode
R4698 N4697 N4698 10
D4698 N4698 0 diode
R4699 N4698 N4699 10
D4699 N4699 0 diode
R4700 N4699 N4700 10
D4700 N4700 0 diode
R4701 N4700 N4701 10
D4701 N4701 0 diode
R4702 N4701 N4702 10
D4702 N4702 0 diode
R4703 N4702 N4703 10
D4703 N4703 0 diode
R4704 N4703 N4704 10
D4704 N4704 0 diode
R4705 N4704 N4705 10
D4705 N4705 0 diode
R4706 N4705 N4706 10
D4706 N4706 0 diode
R4707 N4706 N4707 10
D4707 N4707 0 diode
R4708 N4707 N4708 10
D4708 N4708 0 diode
R4709 N4708 N4709 10
D4709 N4709 0 diode
R4710 N4709 N4710 10
D4710 N4710 0 diode
R4711 N4710 N4711 10
D4711 N4711 0 diode
R4712 N4711 N4712 10
D4712 N4712 0 diode
R4713 N4712 N4713 10
D4713 N4713 0 diode
R4714 N4713 N4714 10
D4714 N4714 0 diode
R4715 N4714 N4715 10
D4715 N4715 0 diode
R4716 N4715 N4716 10
D4716 N4716 0 diode
R4717 N4716 N4717 10
D4717 N4717 0 diode
R4718 N4717 N4718 10
D4718 N4718 0 diode
R4719 N4718 N4719 10
D4719 N4719 0 diode
R4720 N4719 N4720 10
D4720 N4720 0 diode
R4721 N4720 N4721 10
D4721 N4721 0 diode
R4722 N4721 N4722 10
D4722 N4722 0 diode
R4723 N4722 N4723 10
D4723 N4723 0 diode
R4724 N4723 N4724 10
D4724 N4724 0 diode
R4725 N4724 N4725 10
D4725 N4725 0 diode
R4726 N4725 N4726 10
D4726 N4726 0 diode
R4727 N4726 N4727 10
D4727 N4727 0 diode
R4728 N4727 N4728 10
D4728 N4728 0 diode
R4729 N4728 N4729 10
D4729 N4729 0 diode
R4730 N4729 N4730 10
D4730 N4730 0 diode
R4731 N4730 N4731 10
D4731 N4731 0 diode
R4732 N4731 N4732 10
D4732 N4732 0 diode
R4733 N4732 N4733 10
D4733 N4733 0 diode
R4734 N4733 N4734 10
D4734 N4734 0 diode
R4735 N4734 N4735 10
D4735 N4735 0 diode
R4736 N4735 N4736 10
D4736 N4736 0 diode
R4737 N4736 N4737 10
D4737 N4737 0 diode
R4738 N4737 N4738 10
D4738 N4738 0 diode
R4739 N4738 N4739 10
D4739 N4739 0 diode
R4740 N4739 N4740 10
D4740 N4740 0 diode
R4741 N4740 N4741 10
D4741 N4741 0 diode
R4742 N4741 N4742 10
D4742 N4742 0 diode
R4743 N4742 N4743 10
D4743 N4743 0 diode
R4744 N4743 N4744 10
D4744 N4744 0 diode
R4745 N4744 N4745 10
D4745 N4745 0 diode
R4746 N4745 N4746 10
D4746 N4746 0 diode
R4747 N4746 N4747 10
D4747 N4747 0 diode
R4748 N4747 N4748 10
D4748 N4748 0 diode
R4749 N4748 N4749 10
D4749 N4749 0 diode
R4750 N4749 N4750 10
D4750 N4750 0 diode
R4751 N4750 N4751 10
D4751 N4751 0 diode
R4752 N4751 N4752 10
D4752 N4752 0 diode
R4753 N4752 N4753 10
D4753 N4753 0 diode
R4754 N4753 N4754 10
D4754 N4754 0 diode
R4755 N4754 N4755 10
D4755 N4755 0 diode
R4756 N4755 N4756 10
D4756 N4756 0 diode
R4757 N4756 N4757 10
D4757 N4757 0 diode
R4758 N4757 N4758 10
D4758 N4758 0 diode
R4759 N4758 N4759 10
D4759 N4759 0 diode
R4760 N4759 N4760 10
D4760 N4760 0 diode
R4761 N4760 N4761 10
D4761 N4761 0 diode
R4762 N4761 N4762 10
D4762 N4762 0 diode
R4763 N4762 N4763 10
D4763 N4763 0 diode
R4764 N4763 N4764 10
D4764 N4764 0 diode
R4765 N4764 N4765 10
D4765 N4765 0 diode
R4766 N4765 N4766 10
D4766 N4766 0 diode
R4767 N4766 N4767 10
D4767 N4767 0 diode
R4768 N4767 N4768 10
D4768 N4768 0 diode
R4769 N4768 N4769 10
D4769 N4769 0 diode
R4770 N4769 N4770 10
D4770 N4770 0 diode
R4771 N4770 N4771 10
D4771 N4771 0 diode
R4772 N4771 N4772 10
D4772 N4772 0 diode
R4773 N4772 N4773 10
D4773 N4773 0 diode
R4774 N4773 N4774 10
D4774 N4774 0 diode
R4775 N4774 N4775 10
D4775 N4775 0 diode
R4776 N4775 N4776 10
D4776 N4776 0 diode
R4777 N4776 N4777 10
D4777 N4777 0 diode
R4778 N4777 N4778 10
D4778 N4778 0 diode
R4779 N4778 N4779 10
D4779 N4779 0 diode
R4780 N4779 N4780 10
D4780 N4780 0 diode
R4781 N4780 N4781 10
D4781 N4781 0 diode
R4782 N4781 N4782 10
D4782 N4782 0 diode
R4783 N4782 N4783 10
D4783 N4783 0 diode
R4784 N4783 N4784 10
D4784 N4784 0 diode
R4785 N4784 N4785 10
D4785 N4785 0 diode
R4786 N4785 N4786 10
D4786 N4786 0 diode
R4787 N4786 N4787 10
D4787 N4787 0 diode
R4788 N4787 N4788 10
D4788 N4788 0 diode
R4789 N4788 N4789 10
D4789 N4789 0 diode
R4790 N4789 N4790 10
D4790 N4790 0 diode
R4791 N4790 N4791 10
D4791 N4791 0 diode
R4792 N4791 N4792 10
D4792 N4792 0 diode
R4793 N4792 N4793 10
D4793 N4793 0 diode
R4794 N4793 N4794 10
D4794 N4794 0 diode
R4795 N4794 N4795 10
D4795 N4795 0 diode
R4796 N4795 N4796 10
D4796 N4796 0 diode
R4797 N4796 N4797 10
D4797 N4797 0 diode
R4798 N4797 N4798 10
D4798 N4798 0 diode
R4799 N4798 N4799 10
D4799 N4799 0 diode
R4800 N4799 N4800 10
D4800 N4800 0 diode
R4801 N4800 N4801 10
D4801 N4801 0 diode
R4802 N4801 N4802 10
D4802 N4802 0 diode
R4803 N4802 N4803 10
D4803 N4803 0 diode
R4804 N4803 N4804 10
D4804 N4804 0 diode
R4805 N4804 N4805 10
D4805 N4805 0 diode
R4806 N4805 N4806 10
D4806 N4806 0 diode
R4807 N4806 N4807 10
D4807 N4807 0 diode
R4808 N4807 N4808 10
D4808 N4808 0 diode
R4809 N4808 N4809 10
D4809 N4809 0 diode
R4810 N4809 N4810 10
D4810 N4810 0 diode
R4811 N4810 N4811 10
D4811 N4811 0 diode
R4812 N4811 N4812 10
D4812 N4812 0 diode
R4813 N4812 N4813 10
D4813 N4813 0 diode
R4814 N4813 N4814 10
D4814 N4814 0 diode
R4815 N4814 N4815 10
D4815 N4815 0 diode
R4816 N4815 N4816 10
D4816 N4816 0 diode
R4817 N4816 N4817 10
D4817 N4817 0 diode
R4818 N4817 N4818 10
D4818 N4818 0 diode
R4819 N4818 N4819 10
D4819 N4819 0 diode
R4820 N4819 N4820 10
D4820 N4820 0 diode
R4821 N4820 N4821 10
D4821 N4821 0 diode
R4822 N4821 N4822 10
D4822 N4822 0 diode
R4823 N4822 N4823 10
D4823 N4823 0 diode
R4824 N4823 N4824 10
D4824 N4824 0 diode
R4825 N4824 N4825 10
D4825 N4825 0 diode
R4826 N4825 N4826 10
D4826 N4826 0 diode
R4827 N4826 N4827 10
D4827 N4827 0 diode
R4828 N4827 N4828 10
D4828 N4828 0 diode
R4829 N4828 N4829 10
D4829 N4829 0 diode
R4830 N4829 N4830 10
D4830 N4830 0 diode
R4831 N4830 N4831 10
D4831 N4831 0 diode
R4832 N4831 N4832 10
D4832 N4832 0 diode
R4833 N4832 N4833 10
D4833 N4833 0 diode
R4834 N4833 N4834 10
D4834 N4834 0 diode
R4835 N4834 N4835 10
D4835 N4835 0 diode
R4836 N4835 N4836 10
D4836 N4836 0 diode
R4837 N4836 N4837 10
D4837 N4837 0 diode
R4838 N4837 N4838 10
D4838 N4838 0 diode
R4839 N4838 N4839 10
D4839 N4839 0 diode
R4840 N4839 N4840 10
D4840 N4840 0 diode
R4841 N4840 N4841 10
D4841 N4841 0 diode
R4842 N4841 N4842 10
D4842 N4842 0 diode
R4843 N4842 N4843 10
D4843 N4843 0 diode
R4844 N4843 N4844 10
D4844 N4844 0 diode
R4845 N4844 N4845 10
D4845 N4845 0 diode
R4846 N4845 N4846 10
D4846 N4846 0 diode
R4847 N4846 N4847 10
D4847 N4847 0 diode
R4848 N4847 N4848 10
D4848 N4848 0 diode
R4849 N4848 N4849 10
D4849 N4849 0 diode
R4850 N4849 N4850 10
D4850 N4850 0 diode
R4851 N4850 N4851 10
D4851 N4851 0 diode
R4852 N4851 N4852 10
D4852 N4852 0 diode
R4853 N4852 N4853 10
D4853 N4853 0 diode
R4854 N4853 N4854 10
D4854 N4854 0 diode
R4855 N4854 N4855 10
D4855 N4855 0 diode
R4856 N4855 N4856 10
D4856 N4856 0 diode
R4857 N4856 N4857 10
D4857 N4857 0 diode
R4858 N4857 N4858 10
D4858 N4858 0 diode
R4859 N4858 N4859 10
D4859 N4859 0 diode
R4860 N4859 N4860 10
D4860 N4860 0 diode
R4861 N4860 N4861 10
D4861 N4861 0 diode
R4862 N4861 N4862 10
D4862 N4862 0 diode
R4863 N4862 N4863 10
D4863 N4863 0 diode
R4864 N4863 N4864 10
D4864 N4864 0 diode
R4865 N4864 N4865 10
D4865 N4865 0 diode
R4866 N4865 N4866 10
D4866 N4866 0 diode
R4867 N4866 N4867 10
D4867 N4867 0 diode
R4868 N4867 N4868 10
D4868 N4868 0 diode
R4869 N4868 N4869 10
D4869 N4869 0 diode
R4870 N4869 N4870 10
D4870 N4870 0 diode
R4871 N4870 N4871 10
D4871 N4871 0 diode
R4872 N4871 N4872 10
D4872 N4872 0 diode
R4873 N4872 N4873 10
D4873 N4873 0 diode
R4874 N4873 N4874 10
D4874 N4874 0 diode
R4875 N4874 N4875 10
D4875 N4875 0 diode
R4876 N4875 N4876 10
D4876 N4876 0 diode
R4877 N4876 N4877 10
D4877 N4877 0 diode
R4878 N4877 N4878 10
D4878 N4878 0 diode
R4879 N4878 N4879 10
D4879 N4879 0 diode
R4880 N4879 N4880 10
D4880 N4880 0 diode
R4881 N4880 N4881 10
D4881 N4881 0 diode
R4882 N4881 N4882 10
D4882 N4882 0 diode
R4883 N4882 N4883 10
D4883 N4883 0 diode
R4884 N4883 N4884 10
D4884 N4884 0 diode
R4885 N4884 N4885 10
D4885 N4885 0 diode
R4886 N4885 N4886 10
D4886 N4886 0 diode
R4887 N4886 N4887 10
D4887 N4887 0 diode
R4888 N4887 N4888 10
D4888 N4888 0 diode
R4889 N4888 N4889 10
D4889 N4889 0 diode
R4890 N4889 N4890 10
D4890 N4890 0 diode
R4891 N4890 N4891 10
D4891 N4891 0 diode
R4892 N4891 N4892 10
D4892 N4892 0 diode
R4893 N4892 N4893 10
D4893 N4893 0 diode
R4894 N4893 N4894 10
D4894 N4894 0 diode
R4895 N4894 N4895 10
D4895 N4895 0 diode
R4896 N4895 N4896 10
D4896 N4896 0 diode
R4897 N4896 N4897 10
D4897 N4897 0 diode
R4898 N4897 N4898 10
D4898 N4898 0 diode
R4899 N4898 N4899 10
D4899 N4899 0 diode
R4900 N4899 N4900 10
D4900 N4900 0 diode
R4901 N4900 N4901 10
D4901 N4901 0 diode
R4902 N4901 N4902 10
D4902 N4902 0 diode
R4903 N4902 N4903 10
D4903 N4903 0 diode
R4904 N4903 N4904 10
D4904 N4904 0 diode
R4905 N4904 N4905 10
D4905 N4905 0 diode
R4906 N4905 N4906 10
D4906 N4906 0 diode
R4907 N4906 N4907 10
D4907 N4907 0 diode
R4908 N4907 N4908 10
D4908 N4908 0 diode
R4909 N4908 N4909 10
D4909 N4909 0 diode
R4910 N4909 N4910 10
D4910 N4910 0 diode
R4911 N4910 N4911 10
D4911 N4911 0 diode
R4912 N4911 N4912 10
D4912 N4912 0 diode
R4913 N4912 N4913 10
D4913 N4913 0 diode
R4914 N4913 N4914 10
D4914 N4914 0 diode
R4915 N4914 N4915 10
D4915 N4915 0 diode
R4916 N4915 N4916 10
D4916 N4916 0 diode
R4917 N4916 N4917 10
D4917 N4917 0 diode
R4918 N4917 N4918 10
D4918 N4918 0 diode
R4919 N4918 N4919 10
D4919 N4919 0 diode
R4920 N4919 N4920 10
D4920 N4920 0 diode
R4921 N4920 N4921 10
D4921 N4921 0 diode
R4922 N4921 N4922 10
D4922 N4922 0 diode
R4923 N4922 N4923 10
D4923 N4923 0 diode
R4924 N4923 N4924 10
D4924 N4924 0 diode
R4925 N4924 N4925 10
D4925 N4925 0 diode
R4926 N4925 N4926 10
D4926 N4926 0 diode
R4927 N4926 N4927 10
D4927 N4927 0 diode
R4928 N4927 N4928 10
D4928 N4928 0 diode
R4929 N4928 N4929 10
D4929 N4929 0 diode
R4930 N4929 N4930 10
D4930 N4930 0 diode
R4931 N4930 N4931 10
D4931 N4931 0 diode
R4932 N4931 N4932 10
D4932 N4932 0 diode
R4933 N4932 N4933 10
D4933 N4933 0 diode
R4934 N4933 N4934 10
D4934 N4934 0 diode
R4935 N4934 N4935 10
D4935 N4935 0 diode
R4936 N4935 N4936 10
D4936 N4936 0 diode
R4937 N4936 N4937 10
D4937 N4937 0 diode
R4938 N4937 N4938 10
D4938 N4938 0 diode
R4939 N4938 N4939 10
D4939 N4939 0 diode
R4940 N4939 N4940 10
D4940 N4940 0 diode
R4941 N4940 N4941 10
D4941 N4941 0 diode
R4942 N4941 N4942 10
D4942 N4942 0 diode
R4943 N4942 N4943 10
D4943 N4943 0 diode
R4944 N4943 N4944 10
D4944 N4944 0 diode
R4945 N4944 N4945 10
D4945 N4945 0 diode
R4946 N4945 N4946 10
D4946 N4946 0 diode
R4947 N4946 N4947 10
D4947 N4947 0 diode
R4948 N4947 N4948 10
D4948 N4948 0 diode
R4949 N4948 N4949 10
D4949 N4949 0 diode
R4950 N4949 N4950 10
D4950 N4950 0 diode
R4951 N4950 N4951 10
D4951 N4951 0 diode
R4952 N4951 N4952 10
D4952 N4952 0 diode
R4953 N4952 N4953 10
D4953 N4953 0 diode
R4954 N4953 N4954 10
D4954 N4954 0 diode
R4955 N4954 N4955 10
D4955 N4955 0 diode
R4956 N4955 N4956 10
D4956 N4956 0 diode
R4957 N4956 N4957 10
D4957 N4957 0 diode
R4958 N4957 N4958 10
D4958 N4958 0 diode
R4959 N4958 N4959 10
D4959 N4959 0 diode
R4960 N4959 N4960 10
D4960 N4960 0 diode
R4961 N4960 N4961 10
D4961 N4961 0 diode
R4962 N4961 N4962 10
D4962 N4962 0 diode
R4963 N4962 N4963 10
D4963 N4963 0 diode
R4964 N4963 N4964 10
D4964 N4964 0 diode
R4965 N4964 N4965 10
D4965 N4965 0 diode
R4966 N4965 N4966 10
D4966 N4966 0 diode
R4967 N4966 N4967 10
D4967 N4967 0 diode
R4968 N4967 N4968 10
D4968 N4968 0 diode
R4969 N4968 N4969 10
D4969 N4969 0 diode
R4970 N4969 N4970 10
D4970 N4970 0 diode
R4971 N4970 N4971 10
D4971 N4971 0 diode
R4972 N4971 N4972 10
D4972 N4972 0 diode
R4973 N4972 N4973 10
D4973 N4973 0 diode
R4974 N4973 N4974 10
D4974 N4974 0 diode
R4975 N4974 N4975 10
D4975 N4975 0 diode
R4976 N4975 N4976 10
D4976 N4976 0 diode
R4977 N4976 N4977 10
D4977 N4977 0 diode
R4978 N4977 N4978 10
D4978 N4978 0 diode
R4979 N4978 N4979 10
D4979 N4979 0 diode
R4980 N4979 N4980 10
D4980 N4980 0 diode
R4981 N4980 N4981 10
D4981 N4981 0 diode
R4982 N4981 N4982 10
D4982 N4982 0 diode
R4983 N4982 N4983 10
D4983 N4983 0 diode
R4984 N4983 N4984 10
D4984 N4984 0 diode
R4985 N4984 N4985 10
D4985 N4985 0 diode
R4986 N4985 N4986 10
D4986 N4986 0 diode
R4987 N4986 N4987 10
D4987 N4987 0 diode
R4988 N4987 N4988 10
D4988 N4988 0 diode
R4989 N4988 N4989 10
D4989 N4989 0 diode
R4990 N4989 N4990 10
D4990 N4990 0 diode
R4991 N4990 N4991 10
D4991 N4991 0 diode
R4992 N4991 N4992 10
D4992 N4992 0 diode
R4993 N4992 N4993 10
D4993 N4993 0 diode
R4994 N4993 N4994 10
D4994 N4994 0 diode
R4995 N4994 N4995 10
D4995 N4995 0 diode
R4996 N4995 N4996 10
D4996 N4996 0 diode
R4997 N4996 N4997 10
D4997 N4997 0 diode
R4998 N4997 N4998 10
D4998 N4998 0 diode
R4999 N4998 N4999 10
D4999 N4999 0 diode
R5000 N4999 N5000 10
D5000 N5000 0 diode
R5001 N5000 N5001 10
D5001 N5001 0 diode
R5002 N5001 N5002 10
D5002 N5002 0 diode
R5003 N5002 N5003 10
D5003 N5003 0 diode
R5004 N5003 N5004 10
D5004 N5004 0 diode
R5005 N5004 N5005 10
D5005 N5005 0 diode
R5006 N5005 N5006 10
D5006 N5006 0 diode
R5007 N5006 N5007 10
D5007 N5007 0 diode
R5008 N5007 N5008 10
D5008 N5008 0 diode
R5009 N5008 N5009 10
D5009 N5009 0 diode
R5010 N5009 N5010 10
D5010 N5010 0 diode
R5011 N5010 N5011 10
D5011 N5011 0 diode
R5012 N5011 N5012 10
D5012 N5012 0 diode
R5013 N5012 N5013 10
D5013 N5013 0 diode
R5014 N5013 N5014 10
D5014 N5014 0 diode
R5015 N5014 N5015 10
D5015 N5015 0 diode
R5016 N5015 N5016 10
D5016 N5016 0 diode
R5017 N5016 N5017 10
D5017 N5017 0 diode
R5018 N5017 N5018 10
D5018 N5018 0 diode
R5019 N5018 N5019 10
D5019 N5019 0 diode
R5020 N5019 N5020 10
D5020 N5020 0 diode
R5021 N5020 N5021 10
D5021 N5021 0 diode
R5022 N5021 N5022 10
D5022 N5022 0 diode
R5023 N5022 N5023 10
D5023 N5023 0 diode
R5024 N5023 N5024 10
D5024 N5024 0 diode
R5025 N5024 N5025 10
D5025 N5025 0 diode
R5026 N5025 N5026 10
D5026 N5026 0 diode
R5027 N5026 N5027 10
D5027 N5027 0 diode
R5028 N5027 N5028 10
D5028 N5028 0 diode
R5029 N5028 N5029 10
D5029 N5029 0 diode
R5030 N5029 N5030 10
D5030 N5030 0 diode
R5031 N5030 N5031 10
D5031 N5031 0 diode
R5032 N5031 N5032 10
D5032 N5032 0 diode
R5033 N5032 N5033 10
D5033 N5033 0 diode
R5034 N5033 N5034 10
D5034 N5034 0 diode
R5035 N5034 N5035 10
D5035 N5035 0 diode
R5036 N5035 N5036 10
D5036 N5036 0 diode
R5037 N5036 N5037 10
D5037 N5037 0 diode
R5038 N5037 N5038 10
D5038 N5038 0 diode
R5039 N5038 N5039 10
D5039 N5039 0 diode
R5040 N5039 N5040 10
D5040 N5040 0 diode
R5041 N5040 N5041 10
D5041 N5041 0 diode
R5042 N5041 N5042 10
D5042 N5042 0 diode
R5043 N5042 N5043 10
D5043 N5043 0 diode
R5044 N5043 N5044 10
D5044 N5044 0 diode
R5045 N5044 N5045 10
D5045 N5045 0 diode
R5046 N5045 N5046 10
D5046 N5046 0 diode
R5047 N5046 N5047 10
D5047 N5047 0 diode
R5048 N5047 N5048 10
D5048 N5048 0 diode
R5049 N5048 N5049 10
D5049 N5049 0 diode
R5050 N5049 N5050 10
D5050 N5050 0 diode
R5051 N5050 N5051 10
D5051 N5051 0 diode
R5052 N5051 N5052 10
D5052 N5052 0 diode
R5053 N5052 N5053 10
D5053 N5053 0 diode
R5054 N5053 N5054 10
D5054 N5054 0 diode
R5055 N5054 N5055 10
D5055 N5055 0 diode
R5056 N5055 N5056 10
D5056 N5056 0 diode
R5057 N5056 N5057 10
D5057 N5057 0 diode
R5058 N5057 N5058 10
D5058 N5058 0 diode
R5059 N5058 N5059 10
D5059 N5059 0 diode
R5060 N5059 N5060 10
D5060 N5060 0 diode
R5061 N5060 N5061 10
D5061 N5061 0 diode
R5062 N5061 N5062 10
D5062 N5062 0 diode
R5063 N5062 N5063 10
D5063 N5063 0 diode
R5064 N5063 N5064 10
D5064 N5064 0 diode
R5065 N5064 N5065 10
D5065 N5065 0 diode
R5066 N5065 N5066 10
D5066 N5066 0 diode
R5067 N5066 N5067 10
D5067 N5067 0 diode
R5068 N5067 N5068 10
D5068 N5068 0 diode
R5069 N5068 N5069 10
D5069 N5069 0 diode
R5070 N5069 N5070 10
D5070 N5070 0 diode
R5071 N5070 N5071 10
D5071 N5071 0 diode
R5072 N5071 N5072 10
D5072 N5072 0 diode
R5073 N5072 N5073 10
D5073 N5073 0 diode
R5074 N5073 N5074 10
D5074 N5074 0 diode
R5075 N5074 N5075 10
D5075 N5075 0 diode
R5076 N5075 N5076 10
D5076 N5076 0 diode
R5077 N5076 N5077 10
D5077 N5077 0 diode
R5078 N5077 N5078 10
D5078 N5078 0 diode
R5079 N5078 N5079 10
D5079 N5079 0 diode
R5080 N5079 N5080 10
D5080 N5080 0 diode
R5081 N5080 N5081 10
D5081 N5081 0 diode
R5082 N5081 N5082 10
D5082 N5082 0 diode
R5083 N5082 N5083 10
D5083 N5083 0 diode
R5084 N5083 N5084 10
D5084 N5084 0 diode
R5085 N5084 N5085 10
D5085 N5085 0 diode
R5086 N5085 N5086 10
D5086 N5086 0 diode
R5087 N5086 N5087 10
D5087 N5087 0 diode
R5088 N5087 N5088 10
D5088 N5088 0 diode
R5089 N5088 N5089 10
D5089 N5089 0 diode
R5090 N5089 N5090 10
D5090 N5090 0 diode
R5091 N5090 N5091 10
D5091 N5091 0 diode
R5092 N5091 N5092 10
D5092 N5092 0 diode
R5093 N5092 N5093 10
D5093 N5093 0 diode
R5094 N5093 N5094 10
D5094 N5094 0 diode
R5095 N5094 N5095 10
D5095 N5095 0 diode
R5096 N5095 N5096 10
D5096 N5096 0 diode
R5097 N5096 N5097 10
D5097 N5097 0 diode
R5098 N5097 N5098 10
D5098 N5098 0 diode
R5099 N5098 N5099 10
D5099 N5099 0 diode
R5100 N5099 N5100 10
D5100 N5100 0 diode
R5101 N5100 N5101 10
D5101 N5101 0 diode
R5102 N5101 N5102 10
D5102 N5102 0 diode
R5103 N5102 N5103 10
D5103 N5103 0 diode
R5104 N5103 N5104 10
D5104 N5104 0 diode
R5105 N5104 N5105 10
D5105 N5105 0 diode
R5106 N5105 N5106 10
D5106 N5106 0 diode
R5107 N5106 N5107 10
D5107 N5107 0 diode
R5108 N5107 N5108 10
D5108 N5108 0 diode
R5109 N5108 N5109 10
D5109 N5109 0 diode
R5110 N5109 N5110 10
D5110 N5110 0 diode
R5111 N5110 N5111 10
D5111 N5111 0 diode
R5112 N5111 N5112 10
D5112 N5112 0 diode
R5113 N5112 N5113 10
D5113 N5113 0 diode
R5114 N5113 N5114 10
D5114 N5114 0 diode
R5115 N5114 N5115 10
D5115 N5115 0 diode
R5116 N5115 N5116 10
D5116 N5116 0 diode
R5117 N5116 N5117 10
D5117 N5117 0 diode
R5118 N5117 N5118 10
D5118 N5118 0 diode
R5119 N5118 N5119 10
D5119 N5119 0 diode
R5120 N5119 N5120 10
D5120 N5120 0 diode
R5121 N5120 N5121 10
D5121 N5121 0 diode
R5122 N5121 N5122 10
D5122 N5122 0 diode
R5123 N5122 N5123 10
D5123 N5123 0 diode
R5124 N5123 N5124 10
D5124 N5124 0 diode
R5125 N5124 N5125 10
D5125 N5125 0 diode
R5126 N5125 N5126 10
D5126 N5126 0 diode
R5127 N5126 N5127 10
D5127 N5127 0 diode
R5128 N5127 N5128 10
D5128 N5128 0 diode
R5129 N5128 N5129 10
D5129 N5129 0 diode
R5130 N5129 N5130 10
D5130 N5130 0 diode
R5131 N5130 N5131 10
D5131 N5131 0 diode
R5132 N5131 N5132 10
D5132 N5132 0 diode
R5133 N5132 N5133 10
D5133 N5133 0 diode
R5134 N5133 N5134 10
D5134 N5134 0 diode
R5135 N5134 N5135 10
D5135 N5135 0 diode
R5136 N5135 N5136 10
D5136 N5136 0 diode
R5137 N5136 N5137 10
D5137 N5137 0 diode
R5138 N5137 N5138 10
D5138 N5138 0 diode
R5139 N5138 N5139 10
D5139 N5139 0 diode
R5140 N5139 N5140 10
D5140 N5140 0 diode
R5141 N5140 N5141 10
D5141 N5141 0 diode
R5142 N5141 N5142 10
D5142 N5142 0 diode
R5143 N5142 N5143 10
D5143 N5143 0 diode
R5144 N5143 N5144 10
D5144 N5144 0 diode
R5145 N5144 N5145 10
D5145 N5145 0 diode
R5146 N5145 N5146 10
D5146 N5146 0 diode
R5147 N5146 N5147 10
D5147 N5147 0 diode
R5148 N5147 N5148 10
D5148 N5148 0 diode
R5149 N5148 N5149 10
D5149 N5149 0 diode
R5150 N5149 N5150 10
D5150 N5150 0 diode
R5151 N5150 N5151 10
D5151 N5151 0 diode
R5152 N5151 N5152 10
D5152 N5152 0 diode
R5153 N5152 N5153 10
D5153 N5153 0 diode
R5154 N5153 N5154 10
D5154 N5154 0 diode
R5155 N5154 N5155 10
D5155 N5155 0 diode
R5156 N5155 N5156 10
D5156 N5156 0 diode
R5157 N5156 N5157 10
D5157 N5157 0 diode
R5158 N5157 N5158 10
D5158 N5158 0 diode
R5159 N5158 N5159 10
D5159 N5159 0 diode
R5160 N5159 N5160 10
D5160 N5160 0 diode
R5161 N5160 N5161 10
D5161 N5161 0 diode
R5162 N5161 N5162 10
D5162 N5162 0 diode
R5163 N5162 N5163 10
D5163 N5163 0 diode
R5164 N5163 N5164 10
D5164 N5164 0 diode
R5165 N5164 N5165 10
D5165 N5165 0 diode
R5166 N5165 N5166 10
D5166 N5166 0 diode
R5167 N5166 N5167 10
D5167 N5167 0 diode
R5168 N5167 N5168 10
D5168 N5168 0 diode
R5169 N5168 N5169 10
D5169 N5169 0 diode
R5170 N5169 N5170 10
D5170 N5170 0 diode
R5171 N5170 N5171 10
D5171 N5171 0 diode
R5172 N5171 N5172 10
D5172 N5172 0 diode
R5173 N5172 N5173 10
D5173 N5173 0 diode
R5174 N5173 N5174 10
D5174 N5174 0 diode
R5175 N5174 N5175 10
D5175 N5175 0 diode
R5176 N5175 N5176 10
D5176 N5176 0 diode
R5177 N5176 N5177 10
D5177 N5177 0 diode
R5178 N5177 N5178 10
D5178 N5178 0 diode
R5179 N5178 N5179 10
D5179 N5179 0 diode
R5180 N5179 N5180 10
D5180 N5180 0 diode
R5181 N5180 N5181 10
D5181 N5181 0 diode
R5182 N5181 N5182 10
D5182 N5182 0 diode
R5183 N5182 N5183 10
D5183 N5183 0 diode
R5184 N5183 N5184 10
D5184 N5184 0 diode
R5185 N5184 N5185 10
D5185 N5185 0 diode
R5186 N5185 N5186 10
D5186 N5186 0 diode
R5187 N5186 N5187 10
D5187 N5187 0 diode
R5188 N5187 N5188 10
D5188 N5188 0 diode
R5189 N5188 N5189 10
D5189 N5189 0 diode
R5190 N5189 N5190 10
D5190 N5190 0 diode
R5191 N5190 N5191 10
D5191 N5191 0 diode
R5192 N5191 N5192 10
D5192 N5192 0 diode
R5193 N5192 N5193 10
D5193 N5193 0 diode
R5194 N5193 N5194 10
D5194 N5194 0 diode
R5195 N5194 N5195 10
D5195 N5195 0 diode
R5196 N5195 N5196 10
D5196 N5196 0 diode
R5197 N5196 N5197 10
D5197 N5197 0 diode
R5198 N5197 N5198 10
D5198 N5198 0 diode
R5199 N5198 N5199 10
D5199 N5199 0 diode
R5200 N5199 N5200 10
D5200 N5200 0 diode
R5201 N5200 N5201 10
D5201 N5201 0 diode
R5202 N5201 N5202 10
D5202 N5202 0 diode
R5203 N5202 N5203 10
D5203 N5203 0 diode
R5204 N5203 N5204 10
D5204 N5204 0 diode
R5205 N5204 N5205 10
D5205 N5205 0 diode
R5206 N5205 N5206 10
D5206 N5206 0 diode
R5207 N5206 N5207 10
D5207 N5207 0 diode
R5208 N5207 N5208 10
D5208 N5208 0 diode
R5209 N5208 N5209 10
D5209 N5209 0 diode
R5210 N5209 N5210 10
D5210 N5210 0 diode
R5211 N5210 N5211 10
D5211 N5211 0 diode
R5212 N5211 N5212 10
D5212 N5212 0 diode
R5213 N5212 N5213 10
D5213 N5213 0 diode
R5214 N5213 N5214 10
D5214 N5214 0 diode
R5215 N5214 N5215 10
D5215 N5215 0 diode
R5216 N5215 N5216 10
D5216 N5216 0 diode
R5217 N5216 N5217 10
D5217 N5217 0 diode
R5218 N5217 N5218 10
D5218 N5218 0 diode
R5219 N5218 N5219 10
D5219 N5219 0 diode
R5220 N5219 N5220 10
D5220 N5220 0 diode
R5221 N5220 N5221 10
D5221 N5221 0 diode
R5222 N5221 N5222 10
D5222 N5222 0 diode
R5223 N5222 N5223 10
D5223 N5223 0 diode
R5224 N5223 N5224 10
D5224 N5224 0 diode
R5225 N5224 N5225 10
D5225 N5225 0 diode
R5226 N5225 N5226 10
D5226 N5226 0 diode
R5227 N5226 N5227 10
D5227 N5227 0 diode
R5228 N5227 N5228 10
D5228 N5228 0 diode
R5229 N5228 N5229 10
D5229 N5229 0 diode
R5230 N5229 N5230 10
D5230 N5230 0 diode
R5231 N5230 N5231 10
D5231 N5231 0 diode
R5232 N5231 N5232 10
D5232 N5232 0 diode
R5233 N5232 N5233 10
D5233 N5233 0 diode
R5234 N5233 N5234 10
D5234 N5234 0 diode
R5235 N5234 N5235 10
D5235 N5235 0 diode
R5236 N5235 N5236 10
D5236 N5236 0 diode
R5237 N5236 N5237 10
D5237 N5237 0 diode
R5238 N5237 N5238 10
D5238 N5238 0 diode
R5239 N5238 N5239 10
D5239 N5239 0 diode
R5240 N5239 N5240 10
D5240 N5240 0 diode
R5241 N5240 N5241 10
D5241 N5241 0 diode
R5242 N5241 N5242 10
D5242 N5242 0 diode
R5243 N5242 N5243 10
D5243 N5243 0 diode
R5244 N5243 N5244 10
D5244 N5244 0 diode
R5245 N5244 N5245 10
D5245 N5245 0 diode
R5246 N5245 N5246 10
D5246 N5246 0 diode
R5247 N5246 N5247 10
D5247 N5247 0 diode
R5248 N5247 N5248 10
D5248 N5248 0 diode
R5249 N5248 N5249 10
D5249 N5249 0 diode
R5250 N5249 N5250 10
D5250 N5250 0 diode
R5251 N5250 N5251 10
D5251 N5251 0 diode
R5252 N5251 N5252 10
D5252 N5252 0 diode
R5253 N5252 N5253 10
D5253 N5253 0 diode
R5254 N5253 N5254 10
D5254 N5254 0 diode
R5255 N5254 N5255 10
D5255 N5255 0 diode
R5256 N5255 N5256 10
D5256 N5256 0 diode
R5257 N5256 N5257 10
D5257 N5257 0 diode
R5258 N5257 N5258 10
D5258 N5258 0 diode
R5259 N5258 N5259 10
D5259 N5259 0 diode
R5260 N5259 N5260 10
D5260 N5260 0 diode
R5261 N5260 N5261 10
D5261 N5261 0 diode
R5262 N5261 N5262 10
D5262 N5262 0 diode
R5263 N5262 N5263 10
D5263 N5263 0 diode
R5264 N5263 N5264 10
D5264 N5264 0 diode
R5265 N5264 N5265 10
D5265 N5265 0 diode
R5266 N5265 N5266 10
D5266 N5266 0 diode
R5267 N5266 N5267 10
D5267 N5267 0 diode
R5268 N5267 N5268 10
D5268 N5268 0 diode
R5269 N5268 N5269 10
D5269 N5269 0 diode
R5270 N5269 N5270 10
D5270 N5270 0 diode
R5271 N5270 N5271 10
D5271 N5271 0 diode
R5272 N5271 N5272 10
D5272 N5272 0 diode
R5273 N5272 N5273 10
D5273 N5273 0 diode
R5274 N5273 N5274 10
D5274 N5274 0 diode
R5275 N5274 N5275 10
D5275 N5275 0 diode
R5276 N5275 N5276 10
D5276 N5276 0 diode
R5277 N5276 N5277 10
D5277 N5277 0 diode
R5278 N5277 N5278 10
D5278 N5278 0 diode
R5279 N5278 N5279 10
D5279 N5279 0 diode
R5280 N5279 N5280 10
D5280 N5280 0 diode
R5281 N5280 N5281 10
D5281 N5281 0 diode
R5282 N5281 N5282 10
D5282 N5282 0 diode
R5283 N5282 N5283 10
D5283 N5283 0 diode
R5284 N5283 N5284 10
D5284 N5284 0 diode
R5285 N5284 N5285 10
D5285 N5285 0 diode
R5286 N5285 N5286 10
D5286 N5286 0 diode
R5287 N5286 N5287 10
D5287 N5287 0 diode
R5288 N5287 N5288 10
D5288 N5288 0 diode
R5289 N5288 N5289 10
D5289 N5289 0 diode
R5290 N5289 N5290 10
D5290 N5290 0 diode
R5291 N5290 N5291 10
D5291 N5291 0 diode
R5292 N5291 N5292 10
D5292 N5292 0 diode
R5293 N5292 N5293 10
D5293 N5293 0 diode
R5294 N5293 N5294 10
D5294 N5294 0 diode
R5295 N5294 N5295 10
D5295 N5295 0 diode
R5296 N5295 N5296 10
D5296 N5296 0 diode
R5297 N5296 N5297 10
D5297 N5297 0 diode
R5298 N5297 N5298 10
D5298 N5298 0 diode
R5299 N5298 N5299 10
D5299 N5299 0 diode
R5300 N5299 N5300 10
D5300 N5300 0 diode
R5301 N5300 N5301 10
D5301 N5301 0 diode
R5302 N5301 N5302 10
D5302 N5302 0 diode
R5303 N5302 N5303 10
D5303 N5303 0 diode
R5304 N5303 N5304 10
D5304 N5304 0 diode
R5305 N5304 N5305 10
D5305 N5305 0 diode
R5306 N5305 N5306 10
D5306 N5306 0 diode
R5307 N5306 N5307 10
D5307 N5307 0 diode
R5308 N5307 N5308 10
D5308 N5308 0 diode
R5309 N5308 N5309 10
D5309 N5309 0 diode
R5310 N5309 N5310 10
D5310 N5310 0 diode
R5311 N5310 N5311 10
D5311 N5311 0 diode
R5312 N5311 N5312 10
D5312 N5312 0 diode
R5313 N5312 N5313 10
D5313 N5313 0 diode
R5314 N5313 N5314 10
D5314 N5314 0 diode
R5315 N5314 N5315 10
D5315 N5315 0 diode
R5316 N5315 N5316 10
D5316 N5316 0 diode
R5317 N5316 N5317 10
D5317 N5317 0 diode
R5318 N5317 N5318 10
D5318 N5318 0 diode
R5319 N5318 N5319 10
D5319 N5319 0 diode
R5320 N5319 N5320 10
D5320 N5320 0 diode
R5321 N5320 N5321 10
D5321 N5321 0 diode
R5322 N5321 N5322 10
D5322 N5322 0 diode
R5323 N5322 N5323 10
D5323 N5323 0 diode
R5324 N5323 N5324 10
D5324 N5324 0 diode
R5325 N5324 N5325 10
D5325 N5325 0 diode
R5326 N5325 N5326 10
D5326 N5326 0 diode
R5327 N5326 N5327 10
D5327 N5327 0 diode
R5328 N5327 N5328 10
D5328 N5328 0 diode
R5329 N5328 N5329 10
D5329 N5329 0 diode
R5330 N5329 N5330 10
D5330 N5330 0 diode
R5331 N5330 N5331 10
D5331 N5331 0 diode
R5332 N5331 N5332 10
D5332 N5332 0 diode
R5333 N5332 N5333 10
D5333 N5333 0 diode
R5334 N5333 N5334 10
D5334 N5334 0 diode
R5335 N5334 N5335 10
D5335 N5335 0 diode
R5336 N5335 N5336 10
D5336 N5336 0 diode
R5337 N5336 N5337 10
D5337 N5337 0 diode
R5338 N5337 N5338 10
D5338 N5338 0 diode
R5339 N5338 N5339 10
D5339 N5339 0 diode
R5340 N5339 N5340 10
D5340 N5340 0 diode
R5341 N5340 N5341 10
D5341 N5341 0 diode
R5342 N5341 N5342 10
D5342 N5342 0 diode
R5343 N5342 N5343 10
D5343 N5343 0 diode
R5344 N5343 N5344 10
D5344 N5344 0 diode
R5345 N5344 N5345 10
D5345 N5345 0 diode
R5346 N5345 N5346 10
D5346 N5346 0 diode
R5347 N5346 N5347 10
D5347 N5347 0 diode
R5348 N5347 N5348 10
D5348 N5348 0 diode
R5349 N5348 N5349 10
D5349 N5349 0 diode
R5350 N5349 N5350 10
D5350 N5350 0 diode
R5351 N5350 N5351 10
D5351 N5351 0 diode
R5352 N5351 N5352 10
D5352 N5352 0 diode
R5353 N5352 N5353 10
D5353 N5353 0 diode
R5354 N5353 N5354 10
D5354 N5354 0 diode
R5355 N5354 N5355 10
D5355 N5355 0 diode
R5356 N5355 N5356 10
D5356 N5356 0 diode
R5357 N5356 N5357 10
D5357 N5357 0 diode
R5358 N5357 N5358 10
D5358 N5358 0 diode
R5359 N5358 N5359 10
D5359 N5359 0 diode
R5360 N5359 N5360 10
D5360 N5360 0 diode
R5361 N5360 N5361 10
D5361 N5361 0 diode
R5362 N5361 N5362 10
D5362 N5362 0 diode
R5363 N5362 N5363 10
D5363 N5363 0 diode
R5364 N5363 N5364 10
D5364 N5364 0 diode
R5365 N5364 N5365 10
D5365 N5365 0 diode
R5366 N5365 N5366 10
D5366 N5366 0 diode
R5367 N5366 N5367 10
D5367 N5367 0 diode
R5368 N5367 N5368 10
D5368 N5368 0 diode
R5369 N5368 N5369 10
D5369 N5369 0 diode
R5370 N5369 N5370 10
D5370 N5370 0 diode
R5371 N5370 N5371 10
D5371 N5371 0 diode
R5372 N5371 N5372 10
D5372 N5372 0 diode
R5373 N5372 N5373 10
D5373 N5373 0 diode
R5374 N5373 N5374 10
D5374 N5374 0 diode
R5375 N5374 N5375 10
D5375 N5375 0 diode
R5376 N5375 N5376 10
D5376 N5376 0 diode
R5377 N5376 N5377 10
D5377 N5377 0 diode
R5378 N5377 N5378 10
D5378 N5378 0 diode
R5379 N5378 N5379 10
D5379 N5379 0 diode
R5380 N5379 N5380 10
D5380 N5380 0 diode
R5381 N5380 N5381 10
D5381 N5381 0 diode
R5382 N5381 N5382 10
D5382 N5382 0 diode
R5383 N5382 N5383 10
D5383 N5383 0 diode
R5384 N5383 N5384 10
D5384 N5384 0 diode
R5385 N5384 N5385 10
D5385 N5385 0 diode
R5386 N5385 N5386 10
D5386 N5386 0 diode
R5387 N5386 N5387 10
D5387 N5387 0 diode
R5388 N5387 N5388 10
D5388 N5388 0 diode
R5389 N5388 N5389 10
D5389 N5389 0 diode
R5390 N5389 N5390 10
D5390 N5390 0 diode
R5391 N5390 N5391 10
D5391 N5391 0 diode
R5392 N5391 N5392 10
D5392 N5392 0 diode
R5393 N5392 N5393 10
D5393 N5393 0 diode
R5394 N5393 N5394 10
D5394 N5394 0 diode
R5395 N5394 N5395 10
D5395 N5395 0 diode
R5396 N5395 N5396 10
D5396 N5396 0 diode
R5397 N5396 N5397 10
D5397 N5397 0 diode
R5398 N5397 N5398 10
D5398 N5398 0 diode
R5399 N5398 N5399 10
D5399 N5399 0 diode
R5400 N5399 N5400 10
D5400 N5400 0 diode
R5401 N5400 N5401 10
D5401 N5401 0 diode
R5402 N5401 N5402 10
D5402 N5402 0 diode
R5403 N5402 N5403 10
D5403 N5403 0 diode
R5404 N5403 N5404 10
D5404 N5404 0 diode
R5405 N5404 N5405 10
D5405 N5405 0 diode
R5406 N5405 N5406 10
D5406 N5406 0 diode
R5407 N5406 N5407 10
D5407 N5407 0 diode
R5408 N5407 N5408 10
D5408 N5408 0 diode
R5409 N5408 N5409 10
D5409 N5409 0 diode
R5410 N5409 N5410 10
D5410 N5410 0 diode
R5411 N5410 N5411 10
D5411 N5411 0 diode
R5412 N5411 N5412 10
D5412 N5412 0 diode
R5413 N5412 N5413 10
D5413 N5413 0 diode
R5414 N5413 N5414 10
D5414 N5414 0 diode
R5415 N5414 N5415 10
D5415 N5415 0 diode
R5416 N5415 N5416 10
D5416 N5416 0 diode
R5417 N5416 N5417 10
D5417 N5417 0 diode
R5418 N5417 N5418 10
D5418 N5418 0 diode
R5419 N5418 N5419 10
D5419 N5419 0 diode
R5420 N5419 N5420 10
D5420 N5420 0 diode
R5421 N5420 N5421 10
D5421 N5421 0 diode
R5422 N5421 N5422 10
D5422 N5422 0 diode
R5423 N5422 N5423 10
D5423 N5423 0 diode
R5424 N5423 N5424 10
D5424 N5424 0 diode
R5425 N5424 N5425 10
D5425 N5425 0 diode
R5426 N5425 N5426 10
D5426 N5426 0 diode
R5427 N5426 N5427 10
D5427 N5427 0 diode
R5428 N5427 N5428 10
D5428 N5428 0 diode
R5429 N5428 N5429 10
D5429 N5429 0 diode
R5430 N5429 N5430 10
D5430 N5430 0 diode
R5431 N5430 N5431 10
D5431 N5431 0 diode
R5432 N5431 N5432 10
D5432 N5432 0 diode
R5433 N5432 N5433 10
D5433 N5433 0 diode
R5434 N5433 N5434 10
D5434 N5434 0 diode
R5435 N5434 N5435 10
D5435 N5435 0 diode
R5436 N5435 N5436 10
D5436 N5436 0 diode
R5437 N5436 N5437 10
D5437 N5437 0 diode
R5438 N5437 N5438 10
D5438 N5438 0 diode
R5439 N5438 N5439 10
D5439 N5439 0 diode
R5440 N5439 N5440 10
D5440 N5440 0 diode
R5441 N5440 N5441 10
D5441 N5441 0 diode
R5442 N5441 N5442 10
D5442 N5442 0 diode
R5443 N5442 N5443 10
D5443 N5443 0 diode
R5444 N5443 N5444 10
D5444 N5444 0 diode
R5445 N5444 N5445 10
D5445 N5445 0 diode
R5446 N5445 N5446 10
D5446 N5446 0 diode
R5447 N5446 N5447 10
D5447 N5447 0 diode
R5448 N5447 N5448 10
D5448 N5448 0 diode
R5449 N5448 N5449 10
D5449 N5449 0 diode
R5450 N5449 N5450 10
D5450 N5450 0 diode
R5451 N5450 N5451 10
D5451 N5451 0 diode
R5452 N5451 N5452 10
D5452 N5452 0 diode
R5453 N5452 N5453 10
D5453 N5453 0 diode
R5454 N5453 N5454 10
D5454 N5454 0 diode
R5455 N5454 N5455 10
D5455 N5455 0 diode
R5456 N5455 N5456 10
D5456 N5456 0 diode
R5457 N5456 N5457 10
D5457 N5457 0 diode
R5458 N5457 N5458 10
D5458 N5458 0 diode
R5459 N5458 N5459 10
D5459 N5459 0 diode
R5460 N5459 N5460 10
D5460 N5460 0 diode
R5461 N5460 N5461 10
D5461 N5461 0 diode
R5462 N5461 N5462 10
D5462 N5462 0 diode
R5463 N5462 N5463 10
D5463 N5463 0 diode
R5464 N5463 N5464 10
D5464 N5464 0 diode
R5465 N5464 N5465 10
D5465 N5465 0 diode
R5466 N5465 N5466 10
D5466 N5466 0 diode
R5467 N5466 N5467 10
D5467 N5467 0 diode
R5468 N5467 N5468 10
D5468 N5468 0 diode
R5469 N5468 N5469 10
D5469 N5469 0 diode
R5470 N5469 N5470 10
D5470 N5470 0 diode
R5471 N5470 N5471 10
D5471 N5471 0 diode
R5472 N5471 N5472 10
D5472 N5472 0 diode
R5473 N5472 N5473 10
D5473 N5473 0 diode
R5474 N5473 N5474 10
D5474 N5474 0 diode
R5475 N5474 N5475 10
D5475 N5475 0 diode
R5476 N5475 N5476 10
D5476 N5476 0 diode
R5477 N5476 N5477 10
D5477 N5477 0 diode
R5478 N5477 N5478 10
D5478 N5478 0 diode
R5479 N5478 N5479 10
D5479 N5479 0 diode
R5480 N5479 N5480 10
D5480 N5480 0 diode
R5481 N5480 N5481 10
D5481 N5481 0 diode
R5482 N5481 N5482 10
D5482 N5482 0 diode
R5483 N5482 N5483 10
D5483 N5483 0 diode
R5484 N5483 N5484 10
D5484 N5484 0 diode
R5485 N5484 N5485 10
D5485 N5485 0 diode
R5486 N5485 N5486 10
D5486 N5486 0 diode
R5487 N5486 N5487 10
D5487 N5487 0 diode
R5488 N5487 N5488 10
D5488 N5488 0 diode
R5489 N5488 N5489 10
D5489 N5489 0 diode
R5490 N5489 N5490 10
D5490 N5490 0 diode
R5491 N5490 N5491 10
D5491 N5491 0 diode
R5492 N5491 N5492 10
D5492 N5492 0 diode
R5493 N5492 N5493 10
D5493 N5493 0 diode
R5494 N5493 N5494 10
D5494 N5494 0 diode
R5495 N5494 N5495 10
D5495 N5495 0 diode
R5496 N5495 N5496 10
D5496 N5496 0 diode
R5497 N5496 N5497 10
D5497 N5497 0 diode
R5498 N5497 N5498 10
D5498 N5498 0 diode
R5499 N5498 N5499 10
D5499 N5499 0 diode
R5500 N5499 N5500 10
D5500 N5500 0 diode
R5501 N5500 N5501 10
D5501 N5501 0 diode
R5502 N5501 N5502 10
D5502 N5502 0 diode
R5503 N5502 N5503 10
D5503 N5503 0 diode
R5504 N5503 N5504 10
D5504 N5504 0 diode
R5505 N5504 N5505 10
D5505 N5505 0 diode
R5506 N5505 N5506 10
D5506 N5506 0 diode
R5507 N5506 N5507 10
D5507 N5507 0 diode
R5508 N5507 N5508 10
D5508 N5508 0 diode
R5509 N5508 N5509 10
D5509 N5509 0 diode
R5510 N5509 N5510 10
D5510 N5510 0 diode
R5511 N5510 N5511 10
D5511 N5511 0 diode
R5512 N5511 N5512 10
D5512 N5512 0 diode
R5513 N5512 N5513 10
D5513 N5513 0 diode
R5514 N5513 N5514 10
D5514 N5514 0 diode
R5515 N5514 N5515 10
D5515 N5515 0 diode
R5516 N5515 N5516 10
D5516 N5516 0 diode
R5517 N5516 N5517 10
D5517 N5517 0 diode
R5518 N5517 N5518 10
D5518 N5518 0 diode
R5519 N5518 N5519 10
D5519 N5519 0 diode
R5520 N5519 N5520 10
D5520 N5520 0 diode
R5521 N5520 N5521 10
D5521 N5521 0 diode
R5522 N5521 N5522 10
D5522 N5522 0 diode
R5523 N5522 N5523 10
D5523 N5523 0 diode
R5524 N5523 N5524 10
D5524 N5524 0 diode
R5525 N5524 N5525 10
D5525 N5525 0 diode
R5526 N5525 N5526 10
D5526 N5526 0 diode
R5527 N5526 N5527 10
D5527 N5527 0 diode
R5528 N5527 N5528 10
D5528 N5528 0 diode
R5529 N5528 N5529 10
D5529 N5529 0 diode
R5530 N5529 N5530 10
D5530 N5530 0 diode
R5531 N5530 N5531 10
D5531 N5531 0 diode
R5532 N5531 N5532 10
D5532 N5532 0 diode
R5533 N5532 N5533 10
D5533 N5533 0 diode
R5534 N5533 N5534 10
D5534 N5534 0 diode
R5535 N5534 N5535 10
D5535 N5535 0 diode
R5536 N5535 N5536 10
D5536 N5536 0 diode
R5537 N5536 N5537 10
D5537 N5537 0 diode
R5538 N5537 N5538 10
D5538 N5538 0 diode
R5539 N5538 N5539 10
D5539 N5539 0 diode
R5540 N5539 N5540 10
D5540 N5540 0 diode
R5541 N5540 N5541 10
D5541 N5541 0 diode
R5542 N5541 N5542 10
D5542 N5542 0 diode
R5543 N5542 N5543 10
D5543 N5543 0 diode
R5544 N5543 N5544 10
D5544 N5544 0 diode
R5545 N5544 N5545 10
D5545 N5545 0 diode
R5546 N5545 N5546 10
D5546 N5546 0 diode
R5547 N5546 N5547 10
D5547 N5547 0 diode
R5548 N5547 N5548 10
D5548 N5548 0 diode
R5549 N5548 N5549 10
D5549 N5549 0 diode
R5550 N5549 N5550 10
D5550 N5550 0 diode
R5551 N5550 N5551 10
D5551 N5551 0 diode
R5552 N5551 N5552 10
D5552 N5552 0 diode
R5553 N5552 N5553 10
D5553 N5553 0 diode
R5554 N5553 N5554 10
D5554 N5554 0 diode
R5555 N5554 N5555 10
D5555 N5555 0 diode
R5556 N5555 N5556 10
D5556 N5556 0 diode
R5557 N5556 N5557 10
D5557 N5557 0 diode
R5558 N5557 N5558 10
D5558 N5558 0 diode
R5559 N5558 N5559 10
D5559 N5559 0 diode
R5560 N5559 N5560 10
D5560 N5560 0 diode
R5561 N5560 N5561 10
D5561 N5561 0 diode
R5562 N5561 N5562 10
D5562 N5562 0 diode
R5563 N5562 N5563 10
D5563 N5563 0 diode
R5564 N5563 N5564 10
D5564 N5564 0 diode
R5565 N5564 N5565 10
D5565 N5565 0 diode
R5566 N5565 N5566 10
D5566 N5566 0 diode
R5567 N5566 N5567 10
D5567 N5567 0 diode
R5568 N5567 N5568 10
D5568 N5568 0 diode
R5569 N5568 N5569 10
D5569 N5569 0 diode
R5570 N5569 N5570 10
D5570 N5570 0 diode
R5571 N5570 N5571 10
D5571 N5571 0 diode
R5572 N5571 N5572 10
D5572 N5572 0 diode
R5573 N5572 N5573 10
D5573 N5573 0 diode
R5574 N5573 N5574 10
D5574 N5574 0 diode
R5575 N5574 N5575 10
D5575 N5575 0 diode
R5576 N5575 N5576 10
D5576 N5576 0 diode
R5577 N5576 N5577 10
D5577 N5577 0 diode
R5578 N5577 N5578 10
D5578 N5578 0 diode
R5579 N5578 N5579 10
D5579 N5579 0 diode
R5580 N5579 N5580 10
D5580 N5580 0 diode
R5581 N5580 N5581 10
D5581 N5581 0 diode
R5582 N5581 N5582 10
D5582 N5582 0 diode
R5583 N5582 N5583 10
D5583 N5583 0 diode
R5584 N5583 N5584 10
D5584 N5584 0 diode
R5585 N5584 N5585 10
D5585 N5585 0 diode
R5586 N5585 N5586 10
D5586 N5586 0 diode
R5587 N5586 N5587 10
D5587 N5587 0 diode
R5588 N5587 N5588 10
D5588 N5588 0 diode
R5589 N5588 N5589 10
D5589 N5589 0 diode
R5590 N5589 N5590 10
D5590 N5590 0 diode
R5591 N5590 N5591 10
D5591 N5591 0 diode
R5592 N5591 N5592 10
D5592 N5592 0 diode
R5593 N5592 N5593 10
D5593 N5593 0 diode
R5594 N5593 N5594 10
D5594 N5594 0 diode
R5595 N5594 N5595 10
D5595 N5595 0 diode
R5596 N5595 N5596 10
D5596 N5596 0 diode
R5597 N5596 N5597 10
D5597 N5597 0 diode
R5598 N5597 N5598 10
D5598 N5598 0 diode
R5599 N5598 N5599 10
D5599 N5599 0 diode
R5600 N5599 N5600 10
D5600 N5600 0 diode
R5601 N5600 N5601 10
D5601 N5601 0 diode
R5602 N5601 N5602 10
D5602 N5602 0 diode
R5603 N5602 N5603 10
D5603 N5603 0 diode
R5604 N5603 N5604 10
D5604 N5604 0 diode
R5605 N5604 N5605 10
D5605 N5605 0 diode
R5606 N5605 N5606 10
D5606 N5606 0 diode
R5607 N5606 N5607 10
D5607 N5607 0 diode
R5608 N5607 N5608 10
D5608 N5608 0 diode
R5609 N5608 N5609 10
D5609 N5609 0 diode
R5610 N5609 N5610 10
D5610 N5610 0 diode
R5611 N5610 N5611 10
D5611 N5611 0 diode
R5612 N5611 N5612 10
D5612 N5612 0 diode
R5613 N5612 N5613 10
D5613 N5613 0 diode
R5614 N5613 N5614 10
D5614 N5614 0 diode
R5615 N5614 N5615 10
D5615 N5615 0 diode
R5616 N5615 N5616 10
D5616 N5616 0 diode
R5617 N5616 N5617 10
D5617 N5617 0 diode
R5618 N5617 N5618 10
D5618 N5618 0 diode
R5619 N5618 N5619 10
D5619 N5619 0 diode
R5620 N5619 N5620 10
D5620 N5620 0 diode
R5621 N5620 N5621 10
D5621 N5621 0 diode
R5622 N5621 N5622 10
D5622 N5622 0 diode
R5623 N5622 N5623 10
D5623 N5623 0 diode
R5624 N5623 N5624 10
D5624 N5624 0 diode
R5625 N5624 N5625 10
D5625 N5625 0 diode
R5626 N5625 N5626 10
D5626 N5626 0 diode
R5627 N5626 N5627 10
D5627 N5627 0 diode
R5628 N5627 N5628 10
D5628 N5628 0 diode
R5629 N5628 N5629 10
D5629 N5629 0 diode
R5630 N5629 N5630 10
D5630 N5630 0 diode
R5631 N5630 N5631 10
D5631 N5631 0 diode
R5632 N5631 N5632 10
D5632 N5632 0 diode
R5633 N5632 N5633 10
D5633 N5633 0 diode
R5634 N5633 N5634 10
D5634 N5634 0 diode
R5635 N5634 N5635 10
D5635 N5635 0 diode
R5636 N5635 N5636 10
D5636 N5636 0 diode
R5637 N5636 N5637 10
D5637 N5637 0 diode
R5638 N5637 N5638 10
D5638 N5638 0 diode
R5639 N5638 N5639 10
D5639 N5639 0 diode
R5640 N5639 N5640 10
D5640 N5640 0 diode
R5641 N5640 N5641 10
D5641 N5641 0 diode
R5642 N5641 N5642 10
D5642 N5642 0 diode
R5643 N5642 N5643 10
D5643 N5643 0 diode
R5644 N5643 N5644 10
D5644 N5644 0 diode
R5645 N5644 N5645 10
D5645 N5645 0 diode
R5646 N5645 N5646 10
D5646 N5646 0 diode
R5647 N5646 N5647 10
D5647 N5647 0 diode
R5648 N5647 N5648 10
D5648 N5648 0 diode
R5649 N5648 N5649 10
D5649 N5649 0 diode
R5650 N5649 N5650 10
D5650 N5650 0 diode
R5651 N5650 N5651 10
D5651 N5651 0 diode
R5652 N5651 N5652 10
D5652 N5652 0 diode
R5653 N5652 N5653 10
D5653 N5653 0 diode
R5654 N5653 N5654 10
D5654 N5654 0 diode
R5655 N5654 N5655 10
D5655 N5655 0 diode
R5656 N5655 N5656 10
D5656 N5656 0 diode
R5657 N5656 N5657 10
D5657 N5657 0 diode
R5658 N5657 N5658 10
D5658 N5658 0 diode
R5659 N5658 N5659 10
D5659 N5659 0 diode
R5660 N5659 N5660 10
D5660 N5660 0 diode
R5661 N5660 N5661 10
D5661 N5661 0 diode
R5662 N5661 N5662 10
D5662 N5662 0 diode
R5663 N5662 N5663 10
D5663 N5663 0 diode
R5664 N5663 N5664 10
D5664 N5664 0 diode
R5665 N5664 N5665 10
D5665 N5665 0 diode
R5666 N5665 N5666 10
D5666 N5666 0 diode
R5667 N5666 N5667 10
D5667 N5667 0 diode
R5668 N5667 N5668 10
D5668 N5668 0 diode
R5669 N5668 N5669 10
D5669 N5669 0 diode
R5670 N5669 N5670 10
D5670 N5670 0 diode
R5671 N5670 N5671 10
D5671 N5671 0 diode
R5672 N5671 N5672 10
D5672 N5672 0 diode
R5673 N5672 N5673 10
D5673 N5673 0 diode
R5674 N5673 N5674 10
D5674 N5674 0 diode
R5675 N5674 N5675 10
D5675 N5675 0 diode
R5676 N5675 N5676 10
D5676 N5676 0 diode
R5677 N5676 N5677 10
D5677 N5677 0 diode
R5678 N5677 N5678 10
D5678 N5678 0 diode
R5679 N5678 N5679 10
D5679 N5679 0 diode
R5680 N5679 N5680 10
D5680 N5680 0 diode
R5681 N5680 N5681 10
D5681 N5681 0 diode
R5682 N5681 N5682 10
D5682 N5682 0 diode
R5683 N5682 N5683 10
D5683 N5683 0 diode
R5684 N5683 N5684 10
D5684 N5684 0 diode
R5685 N5684 N5685 10
D5685 N5685 0 diode
R5686 N5685 N5686 10
D5686 N5686 0 diode
R5687 N5686 N5687 10
D5687 N5687 0 diode
R5688 N5687 N5688 10
D5688 N5688 0 diode
R5689 N5688 N5689 10
D5689 N5689 0 diode
R5690 N5689 N5690 10
D5690 N5690 0 diode
R5691 N5690 N5691 10
D5691 N5691 0 diode
R5692 N5691 N5692 10
D5692 N5692 0 diode
R5693 N5692 N5693 10
D5693 N5693 0 diode
R5694 N5693 N5694 10
D5694 N5694 0 diode
R5695 N5694 N5695 10
D5695 N5695 0 diode
R5696 N5695 N5696 10
D5696 N5696 0 diode
R5697 N5696 N5697 10
D5697 N5697 0 diode
R5698 N5697 N5698 10
D5698 N5698 0 diode
R5699 N5698 N5699 10
D5699 N5699 0 diode
R5700 N5699 N5700 10
D5700 N5700 0 diode
R5701 N5700 N5701 10
D5701 N5701 0 diode
R5702 N5701 N5702 10
D5702 N5702 0 diode
R5703 N5702 N5703 10
D5703 N5703 0 diode
R5704 N5703 N5704 10
D5704 N5704 0 diode
R5705 N5704 N5705 10
D5705 N5705 0 diode
R5706 N5705 N5706 10
D5706 N5706 0 diode
R5707 N5706 N5707 10
D5707 N5707 0 diode
R5708 N5707 N5708 10
D5708 N5708 0 diode
R5709 N5708 N5709 10
D5709 N5709 0 diode
R5710 N5709 N5710 10
D5710 N5710 0 diode
R5711 N5710 N5711 10
D5711 N5711 0 diode
R5712 N5711 N5712 10
D5712 N5712 0 diode
R5713 N5712 N5713 10
D5713 N5713 0 diode
R5714 N5713 N5714 10
D5714 N5714 0 diode
R5715 N5714 N5715 10
D5715 N5715 0 diode
R5716 N5715 N5716 10
D5716 N5716 0 diode
R5717 N5716 N5717 10
D5717 N5717 0 diode
R5718 N5717 N5718 10
D5718 N5718 0 diode
R5719 N5718 N5719 10
D5719 N5719 0 diode
R5720 N5719 N5720 10
D5720 N5720 0 diode
R5721 N5720 N5721 10
D5721 N5721 0 diode
R5722 N5721 N5722 10
D5722 N5722 0 diode
R5723 N5722 N5723 10
D5723 N5723 0 diode
R5724 N5723 N5724 10
D5724 N5724 0 diode
R5725 N5724 N5725 10
D5725 N5725 0 diode
R5726 N5725 N5726 10
D5726 N5726 0 diode
R5727 N5726 N5727 10
D5727 N5727 0 diode
R5728 N5727 N5728 10
D5728 N5728 0 diode
R5729 N5728 N5729 10
D5729 N5729 0 diode
R5730 N5729 N5730 10
D5730 N5730 0 diode
R5731 N5730 N5731 10
D5731 N5731 0 diode
R5732 N5731 N5732 10
D5732 N5732 0 diode
R5733 N5732 N5733 10
D5733 N5733 0 diode
R5734 N5733 N5734 10
D5734 N5734 0 diode
R5735 N5734 N5735 10
D5735 N5735 0 diode
R5736 N5735 N5736 10
D5736 N5736 0 diode
R5737 N5736 N5737 10
D5737 N5737 0 diode
R5738 N5737 N5738 10
D5738 N5738 0 diode
R5739 N5738 N5739 10
D5739 N5739 0 diode
R5740 N5739 N5740 10
D5740 N5740 0 diode
R5741 N5740 N5741 10
D5741 N5741 0 diode
R5742 N5741 N5742 10
D5742 N5742 0 diode
R5743 N5742 N5743 10
D5743 N5743 0 diode
R5744 N5743 N5744 10
D5744 N5744 0 diode
R5745 N5744 N5745 10
D5745 N5745 0 diode
R5746 N5745 N5746 10
D5746 N5746 0 diode
R5747 N5746 N5747 10
D5747 N5747 0 diode
R5748 N5747 N5748 10
D5748 N5748 0 diode
R5749 N5748 N5749 10
D5749 N5749 0 diode
R5750 N5749 N5750 10
D5750 N5750 0 diode
R5751 N5750 N5751 10
D5751 N5751 0 diode
R5752 N5751 N5752 10
D5752 N5752 0 diode
R5753 N5752 N5753 10
D5753 N5753 0 diode
R5754 N5753 N5754 10
D5754 N5754 0 diode
R5755 N5754 N5755 10
D5755 N5755 0 diode
R5756 N5755 N5756 10
D5756 N5756 0 diode
R5757 N5756 N5757 10
D5757 N5757 0 diode
R5758 N5757 N5758 10
D5758 N5758 0 diode
R5759 N5758 N5759 10
D5759 N5759 0 diode
R5760 N5759 N5760 10
D5760 N5760 0 diode
R5761 N5760 N5761 10
D5761 N5761 0 diode
R5762 N5761 N5762 10
D5762 N5762 0 diode
R5763 N5762 N5763 10
D5763 N5763 0 diode
R5764 N5763 N5764 10
D5764 N5764 0 diode
R5765 N5764 N5765 10
D5765 N5765 0 diode
R5766 N5765 N5766 10
D5766 N5766 0 diode
R5767 N5766 N5767 10
D5767 N5767 0 diode
R5768 N5767 N5768 10
D5768 N5768 0 diode
R5769 N5768 N5769 10
D5769 N5769 0 diode
R5770 N5769 N5770 10
D5770 N5770 0 diode
R5771 N5770 N5771 10
D5771 N5771 0 diode
R5772 N5771 N5772 10
D5772 N5772 0 diode
R5773 N5772 N5773 10
D5773 N5773 0 diode
R5774 N5773 N5774 10
D5774 N5774 0 diode
R5775 N5774 N5775 10
D5775 N5775 0 diode
R5776 N5775 N5776 10
D5776 N5776 0 diode
R5777 N5776 N5777 10
D5777 N5777 0 diode
R5778 N5777 N5778 10
D5778 N5778 0 diode
R5779 N5778 N5779 10
D5779 N5779 0 diode
R5780 N5779 N5780 10
D5780 N5780 0 diode
R5781 N5780 N5781 10
D5781 N5781 0 diode
R5782 N5781 N5782 10
D5782 N5782 0 diode
R5783 N5782 N5783 10
D5783 N5783 0 diode
R5784 N5783 N5784 10
D5784 N5784 0 diode
R5785 N5784 N5785 10
D5785 N5785 0 diode
R5786 N5785 N5786 10
D5786 N5786 0 diode
R5787 N5786 N5787 10
D5787 N5787 0 diode
R5788 N5787 N5788 10
D5788 N5788 0 diode
R5789 N5788 N5789 10
D5789 N5789 0 diode
R5790 N5789 N5790 10
D5790 N5790 0 diode
R5791 N5790 N5791 10
D5791 N5791 0 diode
R5792 N5791 N5792 10
D5792 N5792 0 diode
R5793 N5792 N5793 10
D5793 N5793 0 diode
R5794 N5793 N5794 10
D5794 N5794 0 diode
R5795 N5794 N5795 10
D5795 N5795 0 diode
R5796 N5795 N5796 10
D5796 N5796 0 diode
R5797 N5796 N5797 10
D5797 N5797 0 diode
R5798 N5797 N5798 10
D5798 N5798 0 diode
R5799 N5798 N5799 10
D5799 N5799 0 diode
R5800 N5799 N5800 10
D5800 N5800 0 diode
R5801 N5800 N5801 10
D5801 N5801 0 diode
R5802 N5801 N5802 10
D5802 N5802 0 diode
R5803 N5802 N5803 10
D5803 N5803 0 diode
R5804 N5803 N5804 10
D5804 N5804 0 diode
R5805 N5804 N5805 10
D5805 N5805 0 diode
R5806 N5805 N5806 10
D5806 N5806 0 diode
R5807 N5806 N5807 10
D5807 N5807 0 diode
R5808 N5807 N5808 10
D5808 N5808 0 diode
R5809 N5808 N5809 10
D5809 N5809 0 diode
R5810 N5809 N5810 10
D5810 N5810 0 diode
R5811 N5810 N5811 10
D5811 N5811 0 diode
R5812 N5811 N5812 10
D5812 N5812 0 diode
R5813 N5812 N5813 10
D5813 N5813 0 diode
R5814 N5813 N5814 10
D5814 N5814 0 diode
R5815 N5814 N5815 10
D5815 N5815 0 diode
R5816 N5815 N5816 10
D5816 N5816 0 diode
R5817 N5816 N5817 10
D5817 N5817 0 diode
R5818 N5817 N5818 10
D5818 N5818 0 diode
R5819 N5818 N5819 10
D5819 N5819 0 diode
R5820 N5819 N5820 10
D5820 N5820 0 diode
R5821 N5820 N5821 10
D5821 N5821 0 diode
R5822 N5821 N5822 10
D5822 N5822 0 diode
R5823 N5822 N5823 10
D5823 N5823 0 diode
R5824 N5823 N5824 10
D5824 N5824 0 diode
R5825 N5824 N5825 10
D5825 N5825 0 diode
R5826 N5825 N5826 10
D5826 N5826 0 diode
R5827 N5826 N5827 10
D5827 N5827 0 diode
R5828 N5827 N5828 10
D5828 N5828 0 diode
R5829 N5828 N5829 10
D5829 N5829 0 diode
R5830 N5829 N5830 10
D5830 N5830 0 diode
R5831 N5830 N5831 10
D5831 N5831 0 diode
R5832 N5831 N5832 10
D5832 N5832 0 diode
R5833 N5832 N5833 10
D5833 N5833 0 diode
R5834 N5833 N5834 10
D5834 N5834 0 diode
R5835 N5834 N5835 10
D5835 N5835 0 diode
R5836 N5835 N5836 10
D5836 N5836 0 diode
R5837 N5836 N5837 10
D5837 N5837 0 diode
R5838 N5837 N5838 10
D5838 N5838 0 diode
R5839 N5838 N5839 10
D5839 N5839 0 diode
R5840 N5839 N5840 10
D5840 N5840 0 diode
R5841 N5840 N5841 10
D5841 N5841 0 diode
R5842 N5841 N5842 10
D5842 N5842 0 diode
R5843 N5842 N5843 10
D5843 N5843 0 diode
R5844 N5843 N5844 10
D5844 N5844 0 diode
R5845 N5844 N5845 10
D5845 N5845 0 diode
R5846 N5845 N5846 10
D5846 N5846 0 diode
R5847 N5846 N5847 10
D5847 N5847 0 diode
R5848 N5847 N5848 10
D5848 N5848 0 diode
R5849 N5848 N5849 10
D5849 N5849 0 diode
R5850 N5849 N5850 10
D5850 N5850 0 diode
R5851 N5850 N5851 10
D5851 N5851 0 diode
R5852 N5851 N5852 10
D5852 N5852 0 diode
R5853 N5852 N5853 10
D5853 N5853 0 diode
R5854 N5853 N5854 10
D5854 N5854 0 diode
R5855 N5854 N5855 10
D5855 N5855 0 diode
R5856 N5855 N5856 10
D5856 N5856 0 diode
R5857 N5856 N5857 10
D5857 N5857 0 diode
R5858 N5857 N5858 10
D5858 N5858 0 diode
R5859 N5858 N5859 10
D5859 N5859 0 diode
R5860 N5859 N5860 10
D5860 N5860 0 diode
R5861 N5860 N5861 10
D5861 N5861 0 diode
R5862 N5861 N5862 10
D5862 N5862 0 diode
R5863 N5862 N5863 10
D5863 N5863 0 diode
R5864 N5863 N5864 10
D5864 N5864 0 diode
R5865 N5864 N5865 10
D5865 N5865 0 diode
R5866 N5865 N5866 10
D5866 N5866 0 diode
R5867 N5866 N5867 10
D5867 N5867 0 diode
R5868 N5867 N5868 10
D5868 N5868 0 diode
R5869 N5868 N5869 10
D5869 N5869 0 diode
R5870 N5869 N5870 10
D5870 N5870 0 diode
R5871 N5870 N5871 10
D5871 N5871 0 diode
R5872 N5871 N5872 10
D5872 N5872 0 diode
R5873 N5872 N5873 10
D5873 N5873 0 diode
R5874 N5873 N5874 10
D5874 N5874 0 diode
R5875 N5874 N5875 10
D5875 N5875 0 diode
R5876 N5875 N5876 10
D5876 N5876 0 diode
R5877 N5876 N5877 10
D5877 N5877 0 diode
R5878 N5877 N5878 10
D5878 N5878 0 diode
R5879 N5878 N5879 10
D5879 N5879 0 diode
R5880 N5879 N5880 10
D5880 N5880 0 diode
R5881 N5880 N5881 10
D5881 N5881 0 diode
R5882 N5881 N5882 10
D5882 N5882 0 diode
R5883 N5882 N5883 10
D5883 N5883 0 diode
R5884 N5883 N5884 10
D5884 N5884 0 diode
R5885 N5884 N5885 10
D5885 N5885 0 diode
R5886 N5885 N5886 10
D5886 N5886 0 diode
R5887 N5886 N5887 10
D5887 N5887 0 diode
R5888 N5887 N5888 10
D5888 N5888 0 diode
R5889 N5888 N5889 10
D5889 N5889 0 diode
R5890 N5889 N5890 10
D5890 N5890 0 diode
R5891 N5890 N5891 10
D5891 N5891 0 diode
R5892 N5891 N5892 10
D5892 N5892 0 diode
R5893 N5892 N5893 10
D5893 N5893 0 diode
R5894 N5893 N5894 10
D5894 N5894 0 diode
R5895 N5894 N5895 10
D5895 N5895 0 diode
R5896 N5895 N5896 10
D5896 N5896 0 diode
R5897 N5896 N5897 10
D5897 N5897 0 diode
R5898 N5897 N5898 10
D5898 N5898 0 diode
R5899 N5898 N5899 10
D5899 N5899 0 diode
R5900 N5899 N5900 10
D5900 N5900 0 diode
R5901 N5900 N5901 10
D5901 N5901 0 diode
R5902 N5901 N5902 10
D5902 N5902 0 diode
R5903 N5902 N5903 10
D5903 N5903 0 diode
R5904 N5903 N5904 10
D5904 N5904 0 diode
R5905 N5904 N5905 10
D5905 N5905 0 diode
R5906 N5905 N5906 10
D5906 N5906 0 diode
R5907 N5906 N5907 10
D5907 N5907 0 diode
R5908 N5907 N5908 10
D5908 N5908 0 diode
R5909 N5908 N5909 10
D5909 N5909 0 diode
R5910 N5909 N5910 10
D5910 N5910 0 diode
R5911 N5910 N5911 10
D5911 N5911 0 diode
R5912 N5911 N5912 10
D5912 N5912 0 diode
R5913 N5912 N5913 10
D5913 N5913 0 diode
R5914 N5913 N5914 10
D5914 N5914 0 diode
R5915 N5914 N5915 10
D5915 N5915 0 diode
R5916 N5915 N5916 10
D5916 N5916 0 diode
R5917 N5916 N5917 10
D5917 N5917 0 diode
R5918 N5917 N5918 10
D5918 N5918 0 diode
R5919 N5918 N5919 10
D5919 N5919 0 diode
R5920 N5919 N5920 10
D5920 N5920 0 diode
R5921 N5920 N5921 10
D5921 N5921 0 diode
R5922 N5921 N5922 10
D5922 N5922 0 diode
R5923 N5922 N5923 10
D5923 N5923 0 diode
R5924 N5923 N5924 10
D5924 N5924 0 diode
R5925 N5924 N5925 10
D5925 N5925 0 diode
R5926 N5925 N5926 10
D5926 N5926 0 diode
R5927 N5926 N5927 10
D5927 N5927 0 diode
R5928 N5927 N5928 10
D5928 N5928 0 diode
R5929 N5928 N5929 10
D5929 N5929 0 diode
R5930 N5929 N5930 10
D5930 N5930 0 diode
R5931 N5930 N5931 10
D5931 N5931 0 diode
R5932 N5931 N5932 10
D5932 N5932 0 diode
R5933 N5932 N5933 10
D5933 N5933 0 diode
R5934 N5933 N5934 10
D5934 N5934 0 diode
R5935 N5934 N5935 10
D5935 N5935 0 diode
R5936 N5935 N5936 10
D5936 N5936 0 diode
R5937 N5936 N5937 10
D5937 N5937 0 diode
R5938 N5937 N5938 10
D5938 N5938 0 diode
R5939 N5938 N5939 10
D5939 N5939 0 diode
R5940 N5939 N5940 10
D5940 N5940 0 diode
R5941 N5940 N5941 10
D5941 N5941 0 diode
R5942 N5941 N5942 10
D5942 N5942 0 diode
R5943 N5942 N5943 10
D5943 N5943 0 diode
R5944 N5943 N5944 10
D5944 N5944 0 diode
R5945 N5944 N5945 10
D5945 N5945 0 diode
R5946 N5945 N5946 10
D5946 N5946 0 diode
R5947 N5946 N5947 10
D5947 N5947 0 diode
R5948 N5947 N5948 10
D5948 N5948 0 diode
R5949 N5948 N5949 10
D5949 N5949 0 diode
R5950 N5949 N5950 10
D5950 N5950 0 diode
R5951 N5950 N5951 10
D5951 N5951 0 diode
R5952 N5951 N5952 10
D5952 N5952 0 diode
R5953 N5952 N5953 10
D5953 N5953 0 diode
R5954 N5953 N5954 10
D5954 N5954 0 diode
R5955 N5954 N5955 10
D5955 N5955 0 diode
R5956 N5955 N5956 10
D5956 N5956 0 diode
R5957 N5956 N5957 10
D5957 N5957 0 diode
R5958 N5957 N5958 10
D5958 N5958 0 diode
R5959 N5958 N5959 10
D5959 N5959 0 diode
R5960 N5959 N5960 10
D5960 N5960 0 diode
R5961 N5960 N5961 10
D5961 N5961 0 diode
R5962 N5961 N5962 10
D5962 N5962 0 diode
R5963 N5962 N5963 10
D5963 N5963 0 diode
R5964 N5963 N5964 10
D5964 N5964 0 diode
R5965 N5964 N5965 10
D5965 N5965 0 diode
R5966 N5965 N5966 10
D5966 N5966 0 diode
R5967 N5966 N5967 10
D5967 N5967 0 diode
R5968 N5967 N5968 10
D5968 N5968 0 diode
R5969 N5968 N5969 10
D5969 N5969 0 diode
R5970 N5969 N5970 10
D5970 N5970 0 diode
R5971 N5970 N5971 10
D5971 N5971 0 diode
R5972 N5971 N5972 10
D5972 N5972 0 diode
R5973 N5972 N5973 10
D5973 N5973 0 diode
R5974 N5973 N5974 10
D5974 N5974 0 diode
R5975 N5974 N5975 10
D5975 N5975 0 diode
R5976 N5975 N5976 10
D5976 N5976 0 diode
R5977 N5976 N5977 10
D5977 N5977 0 diode
R5978 N5977 N5978 10
D5978 N5978 0 diode
R5979 N5978 N5979 10
D5979 N5979 0 diode
R5980 N5979 N5980 10
D5980 N5980 0 diode
R5981 N5980 N5981 10
D5981 N5981 0 diode
R5982 N5981 N5982 10
D5982 N5982 0 diode
R5983 N5982 N5983 10
D5983 N5983 0 diode
R5984 N5983 N5984 10
D5984 N5984 0 diode
R5985 N5984 N5985 10
D5985 N5985 0 diode
R5986 N5985 N5986 10
D5986 N5986 0 diode
R5987 N5986 N5987 10
D5987 N5987 0 diode
R5988 N5987 N5988 10
D5988 N5988 0 diode
R5989 N5988 N5989 10
D5989 N5989 0 diode
R5990 N5989 N5990 10
D5990 N5990 0 diode
R5991 N5990 N5991 10
D5991 N5991 0 diode
R5992 N5991 N5992 10
D5992 N5992 0 diode
R5993 N5992 N5993 10
D5993 N5993 0 diode
R5994 N5993 N5994 10
D5994 N5994 0 diode
R5995 N5994 N5995 10
D5995 N5995 0 diode
R5996 N5995 N5996 10
D5996 N5996 0 diode
R5997 N5996 N5997 10
D5997 N5997 0 diode
R5998 N5997 N5998 10
D5998 N5998 0 diode
R5999 N5998 N5999 10
D5999 N5999 0 diode
R6000 N5999 N6000 10
D6000 N6000 0 diode
R6001 N6000 N6001 10
D6001 N6001 0 diode
R6002 N6001 N6002 10
D6002 N6002 0 diode
R6003 N6002 N6003 10
D6003 N6003 0 diode
R6004 N6003 N6004 10
D6004 N6004 0 diode
R6005 N6004 N6005 10
D6005 N6005 0 diode
R6006 N6005 N6006 10
D6006 N6006 0 diode
R6007 N6006 N6007 10
D6007 N6007 0 diode
R6008 N6007 N6008 10
D6008 N6008 0 diode
R6009 N6008 N6009 10
D6009 N6009 0 diode
R6010 N6009 N6010 10
D6010 N6010 0 diode
R6011 N6010 N6011 10
D6011 N6011 0 diode
R6012 N6011 N6012 10
D6012 N6012 0 diode
R6013 N6012 N6013 10
D6013 N6013 0 diode
R6014 N6013 N6014 10
D6014 N6014 0 diode
R6015 N6014 N6015 10
D6015 N6015 0 diode
R6016 N6015 N6016 10
D6016 N6016 0 diode
R6017 N6016 N6017 10
D6017 N6017 0 diode
R6018 N6017 N6018 10
D6018 N6018 0 diode
R6019 N6018 N6019 10
D6019 N6019 0 diode
R6020 N6019 N6020 10
D6020 N6020 0 diode
R6021 N6020 N6021 10
D6021 N6021 0 diode
R6022 N6021 N6022 10
D6022 N6022 0 diode
R6023 N6022 N6023 10
D6023 N6023 0 diode
R6024 N6023 N6024 10
D6024 N6024 0 diode
R6025 N6024 N6025 10
D6025 N6025 0 diode
R6026 N6025 N6026 10
D6026 N6026 0 diode
R6027 N6026 N6027 10
D6027 N6027 0 diode
R6028 N6027 N6028 10
D6028 N6028 0 diode
R6029 N6028 N6029 10
D6029 N6029 0 diode
R6030 N6029 N6030 10
D6030 N6030 0 diode
R6031 N6030 N6031 10
D6031 N6031 0 diode
R6032 N6031 N6032 10
D6032 N6032 0 diode
R6033 N6032 N6033 10
D6033 N6033 0 diode
R6034 N6033 N6034 10
D6034 N6034 0 diode
R6035 N6034 N6035 10
D6035 N6035 0 diode
R6036 N6035 N6036 10
D6036 N6036 0 diode
R6037 N6036 N6037 10
D6037 N6037 0 diode
R6038 N6037 N6038 10
D6038 N6038 0 diode
R6039 N6038 N6039 10
D6039 N6039 0 diode
R6040 N6039 N6040 10
D6040 N6040 0 diode
R6041 N6040 N6041 10
D6041 N6041 0 diode
R6042 N6041 N6042 10
D6042 N6042 0 diode
R6043 N6042 N6043 10
D6043 N6043 0 diode
R6044 N6043 N6044 10
D6044 N6044 0 diode
R6045 N6044 N6045 10
D6045 N6045 0 diode
R6046 N6045 N6046 10
D6046 N6046 0 diode
R6047 N6046 N6047 10
D6047 N6047 0 diode
R6048 N6047 N6048 10
D6048 N6048 0 diode
R6049 N6048 N6049 10
D6049 N6049 0 diode
R6050 N6049 N6050 10
D6050 N6050 0 diode
R6051 N6050 N6051 10
D6051 N6051 0 diode
R6052 N6051 N6052 10
D6052 N6052 0 diode
R6053 N6052 N6053 10
D6053 N6053 0 diode
R6054 N6053 N6054 10
D6054 N6054 0 diode
R6055 N6054 N6055 10
D6055 N6055 0 diode
R6056 N6055 N6056 10
D6056 N6056 0 diode
R6057 N6056 N6057 10
D6057 N6057 0 diode
R6058 N6057 N6058 10
D6058 N6058 0 diode
R6059 N6058 N6059 10
D6059 N6059 0 diode
R6060 N6059 N6060 10
D6060 N6060 0 diode
R6061 N6060 N6061 10
D6061 N6061 0 diode
R6062 N6061 N6062 10
D6062 N6062 0 diode
R6063 N6062 N6063 10
D6063 N6063 0 diode
R6064 N6063 N6064 10
D6064 N6064 0 diode
R6065 N6064 N6065 10
D6065 N6065 0 diode
R6066 N6065 N6066 10
D6066 N6066 0 diode
R6067 N6066 N6067 10
D6067 N6067 0 diode
R6068 N6067 N6068 10
D6068 N6068 0 diode
R6069 N6068 N6069 10
D6069 N6069 0 diode
R6070 N6069 N6070 10
D6070 N6070 0 diode
R6071 N6070 N6071 10
D6071 N6071 0 diode
R6072 N6071 N6072 10
D6072 N6072 0 diode
R6073 N6072 N6073 10
D6073 N6073 0 diode
R6074 N6073 N6074 10
D6074 N6074 0 diode
R6075 N6074 N6075 10
D6075 N6075 0 diode
R6076 N6075 N6076 10
D6076 N6076 0 diode
R6077 N6076 N6077 10
D6077 N6077 0 diode
R6078 N6077 N6078 10
D6078 N6078 0 diode
R6079 N6078 N6079 10
D6079 N6079 0 diode
R6080 N6079 N6080 10
D6080 N6080 0 diode
R6081 N6080 N6081 10
D6081 N6081 0 diode
R6082 N6081 N6082 10
D6082 N6082 0 diode
R6083 N6082 N6083 10
D6083 N6083 0 diode
R6084 N6083 N6084 10
D6084 N6084 0 diode
R6085 N6084 N6085 10
D6085 N6085 0 diode
R6086 N6085 N6086 10
D6086 N6086 0 diode
R6087 N6086 N6087 10
D6087 N6087 0 diode
R6088 N6087 N6088 10
D6088 N6088 0 diode
R6089 N6088 N6089 10
D6089 N6089 0 diode
R6090 N6089 N6090 10
D6090 N6090 0 diode
R6091 N6090 N6091 10
D6091 N6091 0 diode
R6092 N6091 N6092 10
D6092 N6092 0 diode
R6093 N6092 N6093 10
D6093 N6093 0 diode
R6094 N6093 N6094 10
D6094 N6094 0 diode
R6095 N6094 N6095 10
D6095 N6095 0 diode
R6096 N6095 N6096 10
D6096 N6096 0 diode
R6097 N6096 N6097 10
D6097 N6097 0 diode
R6098 N6097 N6098 10
D6098 N6098 0 diode
R6099 N6098 N6099 10
D6099 N6099 0 diode
R6100 N6099 N6100 10
D6100 N6100 0 diode
R6101 N6100 N6101 10
D6101 N6101 0 diode
R6102 N6101 N6102 10
D6102 N6102 0 diode
R6103 N6102 N6103 10
D6103 N6103 0 diode
R6104 N6103 N6104 10
D6104 N6104 0 diode
R6105 N6104 N6105 10
D6105 N6105 0 diode
R6106 N6105 N6106 10
D6106 N6106 0 diode
R6107 N6106 N6107 10
D6107 N6107 0 diode
R6108 N6107 N6108 10
D6108 N6108 0 diode
R6109 N6108 N6109 10
D6109 N6109 0 diode
R6110 N6109 N6110 10
D6110 N6110 0 diode
R6111 N6110 N6111 10
D6111 N6111 0 diode
R6112 N6111 N6112 10
D6112 N6112 0 diode
R6113 N6112 N6113 10
D6113 N6113 0 diode
R6114 N6113 N6114 10
D6114 N6114 0 diode
R6115 N6114 N6115 10
D6115 N6115 0 diode
R6116 N6115 N6116 10
D6116 N6116 0 diode
R6117 N6116 N6117 10
D6117 N6117 0 diode
R6118 N6117 N6118 10
D6118 N6118 0 diode
R6119 N6118 N6119 10
D6119 N6119 0 diode
R6120 N6119 N6120 10
D6120 N6120 0 diode
R6121 N6120 N6121 10
D6121 N6121 0 diode
R6122 N6121 N6122 10
D6122 N6122 0 diode
R6123 N6122 N6123 10
D6123 N6123 0 diode
R6124 N6123 N6124 10
D6124 N6124 0 diode
R6125 N6124 N6125 10
D6125 N6125 0 diode
R6126 N6125 N6126 10
D6126 N6126 0 diode
R6127 N6126 N6127 10
D6127 N6127 0 diode
R6128 N6127 N6128 10
D6128 N6128 0 diode
R6129 N6128 N6129 10
D6129 N6129 0 diode
R6130 N6129 N6130 10
D6130 N6130 0 diode
R6131 N6130 N6131 10
D6131 N6131 0 diode
R6132 N6131 N6132 10
D6132 N6132 0 diode
R6133 N6132 N6133 10
D6133 N6133 0 diode
R6134 N6133 N6134 10
D6134 N6134 0 diode
R6135 N6134 N6135 10
D6135 N6135 0 diode
R6136 N6135 N6136 10
D6136 N6136 0 diode
R6137 N6136 N6137 10
D6137 N6137 0 diode
R6138 N6137 N6138 10
D6138 N6138 0 diode
R6139 N6138 N6139 10
D6139 N6139 0 diode
R6140 N6139 N6140 10
D6140 N6140 0 diode
R6141 N6140 N6141 10
D6141 N6141 0 diode
R6142 N6141 N6142 10
D6142 N6142 0 diode
R6143 N6142 N6143 10
D6143 N6143 0 diode
R6144 N6143 N6144 10
D6144 N6144 0 diode
R6145 N6144 N6145 10
D6145 N6145 0 diode
R6146 N6145 N6146 10
D6146 N6146 0 diode
R6147 N6146 N6147 10
D6147 N6147 0 diode
R6148 N6147 N6148 10
D6148 N6148 0 diode
R6149 N6148 N6149 10
D6149 N6149 0 diode
R6150 N6149 N6150 10
D6150 N6150 0 diode
R6151 N6150 N6151 10
D6151 N6151 0 diode
R6152 N6151 N6152 10
D6152 N6152 0 diode
R6153 N6152 N6153 10
D6153 N6153 0 diode
R6154 N6153 N6154 10
D6154 N6154 0 diode
R6155 N6154 N6155 10
D6155 N6155 0 diode
R6156 N6155 N6156 10
D6156 N6156 0 diode
R6157 N6156 N6157 10
D6157 N6157 0 diode
R6158 N6157 N6158 10
D6158 N6158 0 diode
R6159 N6158 N6159 10
D6159 N6159 0 diode
R6160 N6159 N6160 10
D6160 N6160 0 diode
R6161 N6160 N6161 10
D6161 N6161 0 diode
R6162 N6161 N6162 10
D6162 N6162 0 diode
R6163 N6162 N6163 10
D6163 N6163 0 diode
R6164 N6163 N6164 10
D6164 N6164 0 diode
R6165 N6164 N6165 10
D6165 N6165 0 diode
R6166 N6165 N6166 10
D6166 N6166 0 diode
R6167 N6166 N6167 10
D6167 N6167 0 diode
R6168 N6167 N6168 10
D6168 N6168 0 diode
R6169 N6168 N6169 10
D6169 N6169 0 diode
R6170 N6169 N6170 10
D6170 N6170 0 diode
R6171 N6170 N6171 10
D6171 N6171 0 diode
R6172 N6171 N6172 10
D6172 N6172 0 diode
R6173 N6172 N6173 10
D6173 N6173 0 diode
R6174 N6173 N6174 10
D6174 N6174 0 diode
R6175 N6174 N6175 10
D6175 N6175 0 diode
R6176 N6175 N6176 10
D6176 N6176 0 diode
R6177 N6176 N6177 10
D6177 N6177 0 diode
R6178 N6177 N6178 10
D6178 N6178 0 diode
R6179 N6178 N6179 10
D6179 N6179 0 diode
R6180 N6179 N6180 10
D6180 N6180 0 diode
R6181 N6180 N6181 10
D6181 N6181 0 diode
R6182 N6181 N6182 10
D6182 N6182 0 diode
R6183 N6182 N6183 10
D6183 N6183 0 diode
R6184 N6183 N6184 10
D6184 N6184 0 diode
R6185 N6184 N6185 10
D6185 N6185 0 diode
R6186 N6185 N6186 10
D6186 N6186 0 diode
R6187 N6186 N6187 10
D6187 N6187 0 diode
R6188 N6187 N6188 10
D6188 N6188 0 diode
R6189 N6188 N6189 10
D6189 N6189 0 diode
R6190 N6189 N6190 10
D6190 N6190 0 diode
R6191 N6190 N6191 10
D6191 N6191 0 diode
R6192 N6191 N6192 10
D6192 N6192 0 diode
R6193 N6192 N6193 10
D6193 N6193 0 diode
R6194 N6193 N6194 10
D6194 N6194 0 diode
R6195 N6194 N6195 10
D6195 N6195 0 diode
R6196 N6195 N6196 10
D6196 N6196 0 diode
R6197 N6196 N6197 10
D6197 N6197 0 diode
R6198 N6197 N6198 10
D6198 N6198 0 diode
R6199 N6198 N6199 10
D6199 N6199 0 diode
R6200 N6199 N6200 10
D6200 N6200 0 diode
R6201 N6200 N6201 10
D6201 N6201 0 diode
R6202 N6201 N6202 10
D6202 N6202 0 diode
R6203 N6202 N6203 10
D6203 N6203 0 diode
R6204 N6203 N6204 10
D6204 N6204 0 diode
R6205 N6204 N6205 10
D6205 N6205 0 diode
R6206 N6205 N6206 10
D6206 N6206 0 diode
R6207 N6206 N6207 10
D6207 N6207 0 diode
R6208 N6207 N6208 10
D6208 N6208 0 diode
R6209 N6208 N6209 10
D6209 N6209 0 diode
R6210 N6209 N6210 10
D6210 N6210 0 diode
R6211 N6210 N6211 10
D6211 N6211 0 diode
R6212 N6211 N6212 10
D6212 N6212 0 diode
R6213 N6212 N6213 10
D6213 N6213 0 diode
R6214 N6213 N6214 10
D6214 N6214 0 diode
R6215 N6214 N6215 10
D6215 N6215 0 diode
R6216 N6215 N6216 10
D6216 N6216 0 diode
R6217 N6216 N6217 10
D6217 N6217 0 diode
R6218 N6217 N6218 10
D6218 N6218 0 diode
R6219 N6218 N6219 10
D6219 N6219 0 diode
R6220 N6219 N6220 10
D6220 N6220 0 diode
R6221 N6220 N6221 10
D6221 N6221 0 diode
R6222 N6221 N6222 10
D6222 N6222 0 diode
R6223 N6222 N6223 10
D6223 N6223 0 diode
R6224 N6223 N6224 10
D6224 N6224 0 diode
R6225 N6224 N6225 10
D6225 N6225 0 diode
R6226 N6225 N6226 10
D6226 N6226 0 diode
R6227 N6226 N6227 10
D6227 N6227 0 diode
R6228 N6227 N6228 10
D6228 N6228 0 diode
R6229 N6228 N6229 10
D6229 N6229 0 diode
R6230 N6229 N6230 10
D6230 N6230 0 diode
R6231 N6230 N6231 10
D6231 N6231 0 diode
R6232 N6231 N6232 10
D6232 N6232 0 diode
R6233 N6232 N6233 10
D6233 N6233 0 diode
R6234 N6233 N6234 10
D6234 N6234 0 diode
R6235 N6234 N6235 10
D6235 N6235 0 diode
R6236 N6235 N6236 10
D6236 N6236 0 diode
R6237 N6236 N6237 10
D6237 N6237 0 diode
R6238 N6237 N6238 10
D6238 N6238 0 diode
R6239 N6238 N6239 10
D6239 N6239 0 diode
R6240 N6239 N6240 10
D6240 N6240 0 diode
R6241 N6240 N6241 10
D6241 N6241 0 diode
R6242 N6241 N6242 10
D6242 N6242 0 diode
R6243 N6242 N6243 10
D6243 N6243 0 diode
R6244 N6243 N6244 10
D6244 N6244 0 diode
R6245 N6244 N6245 10
D6245 N6245 0 diode
R6246 N6245 N6246 10
D6246 N6246 0 diode
R6247 N6246 N6247 10
D6247 N6247 0 diode
R6248 N6247 N6248 10
D6248 N6248 0 diode
R6249 N6248 N6249 10
D6249 N6249 0 diode
R6250 N6249 N6250 10
D6250 N6250 0 diode
R6251 N6250 N6251 10
D6251 N6251 0 diode
R6252 N6251 N6252 10
D6252 N6252 0 diode
R6253 N6252 N6253 10
D6253 N6253 0 diode
R6254 N6253 N6254 10
D6254 N6254 0 diode
R6255 N6254 N6255 10
D6255 N6255 0 diode
R6256 N6255 N6256 10
D6256 N6256 0 diode
R6257 N6256 N6257 10
D6257 N6257 0 diode
R6258 N6257 N6258 10
D6258 N6258 0 diode
R6259 N6258 N6259 10
D6259 N6259 0 diode
R6260 N6259 N6260 10
D6260 N6260 0 diode
R6261 N6260 N6261 10
D6261 N6261 0 diode
R6262 N6261 N6262 10
D6262 N6262 0 diode
R6263 N6262 N6263 10
D6263 N6263 0 diode
R6264 N6263 N6264 10
D6264 N6264 0 diode
R6265 N6264 N6265 10
D6265 N6265 0 diode
R6266 N6265 N6266 10
D6266 N6266 0 diode
R6267 N6266 N6267 10
D6267 N6267 0 diode
R6268 N6267 N6268 10
D6268 N6268 0 diode
R6269 N6268 N6269 10
D6269 N6269 0 diode
R6270 N6269 N6270 10
D6270 N6270 0 diode
R6271 N6270 N6271 10
D6271 N6271 0 diode
R6272 N6271 N6272 10
D6272 N6272 0 diode
R6273 N6272 N6273 10
D6273 N6273 0 diode
R6274 N6273 N6274 10
D6274 N6274 0 diode
R6275 N6274 N6275 10
D6275 N6275 0 diode
R6276 N6275 N6276 10
D6276 N6276 0 diode
R6277 N6276 N6277 10
D6277 N6277 0 diode
R6278 N6277 N6278 10
D6278 N6278 0 diode
R6279 N6278 N6279 10
D6279 N6279 0 diode
R6280 N6279 N6280 10
D6280 N6280 0 diode
R6281 N6280 N6281 10
D6281 N6281 0 diode
R6282 N6281 N6282 10
D6282 N6282 0 diode
R6283 N6282 N6283 10
D6283 N6283 0 diode
R6284 N6283 N6284 10
D6284 N6284 0 diode
R6285 N6284 N6285 10
D6285 N6285 0 diode
R6286 N6285 N6286 10
D6286 N6286 0 diode
R6287 N6286 N6287 10
D6287 N6287 0 diode
R6288 N6287 N6288 10
D6288 N6288 0 diode
R6289 N6288 N6289 10
D6289 N6289 0 diode
R6290 N6289 N6290 10
D6290 N6290 0 diode
R6291 N6290 N6291 10
D6291 N6291 0 diode
R6292 N6291 N6292 10
D6292 N6292 0 diode
R6293 N6292 N6293 10
D6293 N6293 0 diode
R6294 N6293 N6294 10
D6294 N6294 0 diode
R6295 N6294 N6295 10
D6295 N6295 0 diode
R6296 N6295 N6296 10
D6296 N6296 0 diode
R6297 N6296 N6297 10
D6297 N6297 0 diode
R6298 N6297 N6298 10
D6298 N6298 0 diode
R6299 N6298 N6299 10
D6299 N6299 0 diode
R6300 N6299 N6300 10
D6300 N6300 0 diode
R6301 N6300 N6301 10
D6301 N6301 0 diode
R6302 N6301 N6302 10
D6302 N6302 0 diode
R6303 N6302 N6303 10
D6303 N6303 0 diode
R6304 N6303 N6304 10
D6304 N6304 0 diode
R6305 N6304 N6305 10
D6305 N6305 0 diode
R6306 N6305 N6306 10
D6306 N6306 0 diode
R6307 N6306 N6307 10
D6307 N6307 0 diode
R6308 N6307 N6308 10
D6308 N6308 0 diode
R6309 N6308 N6309 10
D6309 N6309 0 diode
R6310 N6309 N6310 10
D6310 N6310 0 diode
R6311 N6310 N6311 10
D6311 N6311 0 diode
R6312 N6311 N6312 10
D6312 N6312 0 diode
R6313 N6312 N6313 10
D6313 N6313 0 diode
R6314 N6313 N6314 10
D6314 N6314 0 diode
R6315 N6314 N6315 10
D6315 N6315 0 diode
R6316 N6315 N6316 10
D6316 N6316 0 diode
R6317 N6316 N6317 10
D6317 N6317 0 diode
R6318 N6317 N6318 10
D6318 N6318 0 diode
R6319 N6318 N6319 10
D6319 N6319 0 diode
R6320 N6319 N6320 10
D6320 N6320 0 diode
R6321 N6320 N6321 10
D6321 N6321 0 diode
R6322 N6321 N6322 10
D6322 N6322 0 diode
R6323 N6322 N6323 10
D6323 N6323 0 diode
R6324 N6323 N6324 10
D6324 N6324 0 diode
R6325 N6324 N6325 10
D6325 N6325 0 diode
R6326 N6325 N6326 10
D6326 N6326 0 diode
R6327 N6326 N6327 10
D6327 N6327 0 diode
R6328 N6327 N6328 10
D6328 N6328 0 diode
R6329 N6328 N6329 10
D6329 N6329 0 diode
R6330 N6329 N6330 10
D6330 N6330 0 diode
R6331 N6330 N6331 10
D6331 N6331 0 diode
R6332 N6331 N6332 10
D6332 N6332 0 diode
R6333 N6332 N6333 10
D6333 N6333 0 diode
R6334 N6333 N6334 10
D6334 N6334 0 diode
R6335 N6334 N6335 10
D6335 N6335 0 diode
R6336 N6335 N6336 10
D6336 N6336 0 diode
R6337 N6336 N6337 10
D6337 N6337 0 diode
R6338 N6337 N6338 10
D6338 N6338 0 diode
R6339 N6338 N6339 10
D6339 N6339 0 diode
R6340 N6339 N6340 10
D6340 N6340 0 diode
R6341 N6340 N6341 10
D6341 N6341 0 diode
R6342 N6341 N6342 10
D6342 N6342 0 diode
R6343 N6342 N6343 10
D6343 N6343 0 diode
R6344 N6343 N6344 10
D6344 N6344 0 diode
R6345 N6344 N6345 10
D6345 N6345 0 diode
R6346 N6345 N6346 10
D6346 N6346 0 diode
R6347 N6346 N6347 10
D6347 N6347 0 diode
R6348 N6347 N6348 10
D6348 N6348 0 diode
R6349 N6348 N6349 10
D6349 N6349 0 diode
R6350 N6349 N6350 10
D6350 N6350 0 diode
R6351 N6350 N6351 10
D6351 N6351 0 diode
R6352 N6351 N6352 10
D6352 N6352 0 diode
R6353 N6352 N6353 10
D6353 N6353 0 diode
R6354 N6353 N6354 10
D6354 N6354 0 diode
R6355 N6354 N6355 10
D6355 N6355 0 diode
R6356 N6355 N6356 10
D6356 N6356 0 diode
R6357 N6356 N6357 10
D6357 N6357 0 diode
R6358 N6357 N6358 10
D6358 N6358 0 diode
R6359 N6358 N6359 10
D6359 N6359 0 diode
R6360 N6359 N6360 10
D6360 N6360 0 diode
R6361 N6360 N6361 10
D6361 N6361 0 diode
R6362 N6361 N6362 10
D6362 N6362 0 diode
R6363 N6362 N6363 10
D6363 N6363 0 diode
R6364 N6363 N6364 10
D6364 N6364 0 diode
R6365 N6364 N6365 10
D6365 N6365 0 diode
R6366 N6365 N6366 10
D6366 N6366 0 diode
R6367 N6366 N6367 10
D6367 N6367 0 diode
R6368 N6367 N6368 10
D6368 N6368 0 diode
R6369 N6368 N6369 10
D6369 N6369 0 diode
R6370 N6369 N6370 10
D6370 N6370 0 diode
R6371 N6370 N6371 10
D6371 N6371 0 diode
R6372 N6371 N6372 10
D6372 N6372 0 diode
R6373 N6372 N6373 10
D6373 N6373 0 diode
R6374 N6373 N6374 10
D6374 N6374 0 diode
R6375 N6374 N6375 10
D6375 N6375 0 diode
R6376 N6375 N6376 10
D6376 N6376 0 diode
R6377 N6376 N6377 10
D6377 N6377 0 diode
R6378 N6377 N6378 10
D6378 N6378 0 diode
R6379 N6378 N6379 10
D6379 N6379 0 diode
R6380 N6379 N6380 10
D6380 N6380 0 diode
R6381 N6380 N6381 10
D6381 N6381 0 diode
R6382 N6381 N6382 10
D6382 N6382 0 diode
R6383 N6382 N6383 10
D6383 N6383 0 diode
R6384 N6383 N6384 10
D6384 N6384 0 diode
R6385 N6384 N6385 10
D6385 N6385 0 diode
R6386 N6385 N6386 10
D6386 N6386 0 diode
R6387 N6386 N6387 10
D6387 N6387 0 diode
R6388 N6387 N6388 10
D6388 N6388 0 diode
R6389 N6388 N6389 10
D6389 N6389 0 diode
R6390 N6389 N6390 10
D6390 N6390 0 diode
R6391 N6390 N6391 10
D6391 N6391 0 diode
R6392 N6391 N6392 10
D6392 N6392 0 diode
R6393 N6392 N6393 10
D6393 N6393 0 diode
R6394 N6393 N6394 10
D6394 N6394 0 diode
R6395 N6394 N6395 10
D6395 N6395 0 diode
R6396 N6395 N6396 10
D6396 N6396 0 diode
R6397 N6396 N6397 10
D6397 N6397 0 diode
R6398 N6397 N6398 10
D6398 N6398 0 diode
R6399 N6398 N6399 10
D6399 N6399 0 diode
R6400 N6399 N6400 10
D6400 N6400 0 diode
R6401 N6400 N6401 10
D6401 N6401 0 diode
R6402 N6401 N6402 10
D6402 N6402 0 diode
R6403 N6402 N6403 10
D6403 N6403 0 diode
R6404 N6403 N6404 10
D6404 N6404 0 diode
R6405 N6404 N6405 10
D6405 N6405 0 diode
R6406 N6405 N6406 10
D6406 N6406 0 diode
R6407 N6406 N6407 10
D6407 N6407 0 diode
R6408 N6407 N6408 10
D6408 N6408 0 diode
R6409 N6408 N6409 10
D6409 N6409 0 diode
R6410 N6409 N6410 10
D6410 N6410 0 diode
R6411 N6410 N6411 10
D6411 N6411 0 diode
R6412 N6411 N6412 10
D6412 N6412 0 diode
R6413 N6412 N6413 10
D6413 N6413 0 diode
R6414 N6413 N6414 10
D6414 N6414 0 diode
R6415 N6414 N6415 10
D6415 N6415 0 diode
R6416 N6415 N6416 10
D6416 N6416 0 diode
R6417 N6416 N6417 10
D6417 N6417 0 diode
R6418 N6417 N6418 10
D6418 N6418 0 diode
R6419 N6418 N6419 10
D6419 N6419 0 diode
R6420 N6419 N6420 10
D6420 N6420 0 diode
R6421 N6420 N6421 10
D6421 N6421 0 diode
R6422 N6421 N6422 10
D6422 N6422 0 diode
R6423 N6422 N6423 10
D6423 N6423 0 diode
R6424 N6423 N6424 10
D6424 N6424 0 diode
R6425 N6424 N6425 10
D6425 N6425 0 diode
R6426 N6425 N6426 10
D6426 N6426 0 diode
R6427 N6426 N6427 10
D6427 N6427 0 diode
R6428 N6427 N6428 10
D6428 N6428 0 diode
R6429 N6428 N6429 10
D6429 N6429 0 diode
R6430 N6429 N6430 10
D6430 N6430 0 diode
R6431 N6430 N6431 10
D6431 N6431 0 diode
R6432 N6431 N6432 10
D6432 N6432 0 diode
R6433 N6432 N6433 10
D6433 N6433 0 diode
R6434 N6433 N6434 10
D6434 N6434 0 diode
R6435 N6434 N6435 10
D6435 N6435 0 diode
R6436 N6435 N6436 10
D6436 N6436 0 diode
R6437 N6436 N6437 10
D6437 N6437 0 diode
R6438 N6437 N6438 10
D6438 N6438 0 diode
R6439 N6438 N6439 10
D6439 N6439 0 diode
R6440 N6439 N6440 10
D6440 N6440 0 diode
R6441 N6440 N6441 10
D6441 N6441 0 diode
R6442 N6441 N6442 10
D6442 N6442 0 diode
R6443 N6442 N6443 10
D6443 N6443 0 diode
R6444 N6443 N6444 10
D6444 N6444 0 diode
R6445 N6444 N6445 10
D6445 N6445 0 diode
R6446 N6445 N6446 10
D6446 N6446 0 diode
R6447 N6446 N6447 10
D6447 N6447 0 diode
R6448 N6447 N6448 10
D6448 N6448 0 diode
R6449 N6448 N6449 10
D6449 N6449 0 diode
R6450 N6449 N6450 10
D6450 N6450 0 diode
R6451 N6450 N6451 10
D6451 N6451 0 diode
R6452 N6451 N6452 10
D6452 N6452 0 diode
R6453 N6452 N6453 10
D6453 N6453 0 diode
R6454 N6453 N6454 10
D6454 N6454 0 diode
R6455 N6454 N6455 10
D6455 N6455 0 diode
R6456 N6455 N6456 10
D6456 N6456 0 diode
R6457 N6456 N6457 10
D6457 N6457 0 diode
R6458 N6457 N6458 10
D6458 N6458 0 diode
R6459 N6458 N6459 10
D6459 N6459 0 diode
R6460 N6459 N6460 10
D6460 N6460 0 diode
R6461 N6460 N6461 10
D6461 N6461 0 diode
R6462 N6461 N6462 10
D6462 N6462 0 diode
R6463 N6462 N6463 10
D6463 N6463 0 diode
R6464 N6463 N6464 10
D6464 N6464 0 diode
R6465 N6464 N6465 10
D6465 N6465 0 diode
R6466 N6465 N6466 10
D6466 N6466 0 diode
R6467 N6466 N6467 10
D6467 N6467 0 diode
R6468 N6467 N6468 10
D6468 N6468 0 diode
R6469 N6468 N6469 10
D6469 N6469 0 diode
R6470 N6469 N6470 10
D6470 N6470 0 diode
R6471 N6470 N6471 10
D6471 N6471 0 diode
R6472 N6471 N6472 10
D6472 N6472 0 diode
R6473 N6472 N6473 10
D6473 N6473 0 diode
R6474 N6473 N6474 10
D6474 N6474 0 diode
R6475 N6474 N6475 10
D6475 N6475 0 diode
R6476 N6475 N6476 10
D6476 N6476 0 diode
R6477 N6476 N6477 10
D6477 N6477 0 diode
R6478 N6477 N6478 10
D6478 N6478 0 diode
R6479 N6478 N6479 10
D6479 N6479 0 diode
R6480 N6479 N6480 10
D6480 N6480 0 diode
R6481 N6480 N6481 10
D6481 N6481 0 diode
R6482 N6481 N6482 10
D6482 N6482 0 diode
R6483 N6482 N6483 10
D6483 N6483 0 diode
R6484 N6483 N6484 10
D6484 N6484 0 diode
R6485 N6484 N6485 10
D6485 N6485 0 diode
R6486 N6485 N6486 10
D6486 N6486 0 diode
R6487 N6486 N6487 10
D6487 N6487 0 diode
R6488 N6487 N6488 10
D6488 N6488 0 diode
R6489 N6488 N6489 10
D6489 N6489 0 diode
R6490 N6489 N6490 10
D6490 N6490 0 diode
R6491 N6490 N6491 10
D6491 N6491 0 diode
R6492 N6491 N6492 10
D6492 N6492 0 diode
R6493 N6492 N6493 10
D6493 N6493 0 diode
R6494 N6493 N6494 10
D6494 N6494 0 diode
R6495 N6494 N6495 10
D6495 N6495 0 diode
R6496 N6495 N6496 10
D6496 N6496 0 diode
R6497 N6496 N6497 10
D6497 N6497 0 diode
R6498 N6497 N6498 10
D6498 N6498 0 diode
R6499 N6498 N6499 10
D6499 N6499 0 diode
R6500 N6499 N6500 10
D6500 N6500 0 diode
R6501 N6500 N6501 10
D6501 N6501 0 diode
R6502 N6501 N6502 10
D6502 N6502 0 diode
R6503 N6502 N6503 10
D6503 N6503 0 diode
R6504 N6503 N6504 10
D6504 N6504 0 diode
R6505 N6504 N6505 10
D6505 N6505 0 diode
R6506 N6505 N6506 10
D6506 N6506 0 diode
R6507 N6506 N6507 10
D6507 N6507 0 diode
R6508 N6507 N6508 10
D6508 N6508 0 diode
R6509 N6508 N6509 10
D6509 N6509 0 diode
R6510 N6509 N6510 10
D6510 N6510 0 diode
R6511 N6510 N6511 10
D6511 N6511 0 diode
R6512 N6511 N6512 10
D6512 N6512 0 diode
R6513 N6512 N6513 10
D6513 N6513 0 diode
R6514 N6513 N6514 10
D6514 N6514 0 diode
R6515 N6514 N6515 10
D6515 N6515 0 diode
R6516 N6515 N6516 10
D6516 N6516 0 diode
R6517 N6516 N6517 10
D6517 N6517 0 diode
R6518 N6517 N6518 10
D6518 N6518 0 diode
R6519 N6518 N6519 10
D6519 N6519 0 diode
R6520 N6519 N6520 10
D6520 N6520 0 diode
R6521 N6520 N6521 10
D6521 N6521 0 diode
R6522 N6521 N6522 10
D6522 N6522 0 diode
R6523 N6522 N6523 10
D6523 N6523 0 diode
R6524 N6523 N6524 10
D6524 N6524 0 diode
R6525 N6524 N6525 10
D6525 N6525 0 diode
R6526 N6525 N6526 10
D6526 N6526 0 diode
R6527 N6526 N6527 10
D6527 N6527 0 diode
R6528 N6527 N6528 10
D6528 N6528 0 diode
R6529 N6528 N6529 10
D6529 N6529 0 diode
R6530 N6529 N6530 10
D6530 N6530 0 diode
R6531 N6530 N6531 10
D6531 N6531 0 diode
R6532 N6531 N6532 10
D6532 N6532 0 diode
R6533 N6532 N6533 10
D6533 N6533 0 diode
R6534 N6533 N6534 10
D6534 N6534 0 diode
R6535 N6534 N6535 10
D6535 N6535 0 diode
R6536 N6535 N6536 10
D6536 N6536 0 diode
R6537 N6536 N6537 10
D6537 N6537 0 diode
R6538 N6537 N6538 10
D6538 N6538 0 diode
R6539 N6538 N6539 10
D6539 N6539 0 diode
R6540 N6539 N6540 10
D6540 N6540 0 diode
R6541 N6540 N6541 10
D6541 N6541 0 diode
R6542 N6541 N6542 10
D6542 N6542 0 diode
R6543 N6542 N6543 10
D6543 N6543 0 diode
R6544 N6543 N6544 10
D6544 N6544 0 diode
R6545 N6544 N6545 10
D6545 N6545 0 diode
R6546 N6545 N6546 10
D6546 N6546 0 diode
R6547 N6546 N6547 10
D6547 N6547 0 diode
R6548 N6547 N6548 10
D6548 N6548 0 diode
R6549 N6548 N6549 10
D6549 N6549 0 diode
R6550 N6549 N6550 10
D6550 N6550 0 diode
R6551 N6550 N6551 10
D6551 N6551 0 diode
R6552 N6551 N6552 10
D6552 N6552 0 diode
R6553 N6552 N6553 10
D6553 N6553 0 diode
R6554 N6553 N6554 10
D6554 N6554 0 diode
R6555 N6554 N6555 10
D6555 N6555 0 diode
R6556 N6555 N6556 10
D6556 N6556 0 diode
R6557 N6556 N6557 10
D6557 N6557 0 diode
R6558 N6557 N6558 10
D6558 N6558 0 diode
R6559 N6558 N6559 10
D6559 N6559 0 diode
R6560 N6559 N6560 10
D6560 N6560 0 diode
R6561 N6560 N6561 10
D6561 N6561 0 diode
R6562 N6561 N6562 10
D6562 N6562 0 diode
R6563 N6562 N6563 10
D6563 N6563 0 diode
R6564 N6563 N6564 10
D6564 N6564 0 diode
R6565 N6564 N6565 10
D6565 N6565 0 diode
R6566 N6565 N6566 10
D6566 N6566 0 diode
R6567 N6566 N6567 10
D6567 N6567 0 diode
R6568 N6567 N6568 10
D6568 N6568 0 diode
R6569 N6568 N6569 10
D6569 N6569 0 diode
R6570 N6569 N6570 10
D6570 N6570 0 diode
R6571 N6570 N6571 10
D6571 N6571 0 diode
R6572 N6571 N6572 10
D6572 N6572 0 diode
R6573 N6572 N6573 10
D6573 N6573 0 diode
R6574 N6573 N6574 10
D6574 N6574 0 diode
R6575 N6574 N6575 10
D6575 N6575 0 diode
R6576 N6575 N6576 10
D6576 N6576 0 diode
R6577 N6576 N6577 10
D6577 N6577 0 diode
R6578 N6577 N6578 10
D6578 N6578 0 diode
R6579 N6578 N6579 10
D6579 N6579 0 diode
R6580 N6579 N6580 10
D6580 N6580 0 diode
R6581 N6580 N6581 10
D6581 N6581 0 diode
R6582 N6581 N6582 10
D6582 N6582 0 diode
R6583 N6582 N6583 10
D6583 N6583 0 diode
R6584 N6583 N6584 10
D6584 N6584 0 diode
R6585 N6584 N6585 10
D6585 N6585 0 diode
R6586 N6585 N6586 10
D6586 N6586 0 diode
R6587 N6586 N6587 10
D6587 N6587 0 diode
R6588 N6587 N6588 10
D6588 N6588 0 diode
R6589 N6588 N6589 10
D6589 N6589 0 diode
R6590 N6589 N6590 10
D6590 N6590 0 diode
R6591 N6590 N6591 10
D6591 N6591 0 diode
R6592 N6591 N6592 10
D6592 N6592 0 diode
R6593 N6592 N6593 10
D6593 N6593 0 diode
R6594 N6593 N6594 10
D6594 N6594 0 diode
R6595 N6594 N6595 10
D6595 N6595 0 diode
R6596 N6595 N6596 10
D6596 N6596 0 diode
R6597 N6596 N6597 10
D6597 N6597 0 diode
R6598 N6597 N6598 10
D6598 N6598 0 diode
R6599 N6598 N6599 10
D6599 N6599 0 diode
R6600 N6599 N6600 10
D6600 N6600 0 diode
R6601 N6600 N6601 10
D6601 N6601 0 diode
R6602 N6601 N6602 10
D6602 N6602 0 diode
R6603 N6602 N6603 10
D6603 N6603 0 diode
R6604 N6603 N6604 10
D6604 N6604 0 diode
R6605 N6604 N6605 10
D6605 N6605 0 diode
R6606 N6605 N6606 10
D6606 N6606 0 diode
R6607 N6606 N6607 10
D6607 N6607 0 diode
R6608 N6607 N6608 10
D6608 N6608 0 diode
R6609 N6608 N6609 10
D6609 N6609 0 diode
R6610 N6609 N6610 10
D6610 N6610 0 diode
R6611 N6610 N6611 10
D6611 N6611 0 diode
R6612 N6611 N6612 10
D6612 N6612 0 diode
R6613 N6612 N6613 10
D6613 N6613 0 diode
R6614 N6613 N6614 10
D6614 N6614 0 diode
R6615 N6614 N6615 10
D6615 N6615 0 diode
R6616 N6615 N6616 10
D6616 N6616 0 diode
R6617 N6616 N6617 10
D6617 N6617 0 diode
R6618 N6617 N6618 10
D6618 N6618 0 diode
R6619 N6618 N6619 10
D6619 N6619 0 diode
R6620 N6619 N6620 10
D6620 N6620 0 diode
R6621 N6620 N6621 10
D6621 N6621 0 diode
R6622 N6621 N6622 10
D6622 N6622 0 diode
R6623 N6622 N6623 10
D6623 N6623 0 diode
R6624 N6623 N6624 10
D6624 N6624 0 diode
R6625 N6624 N6625 10
D6625 N6625 0 diode
R6626 N6625 N6626 10
D6626 N6626 0 diode
R6627 N6626 N6627 10
D6627 N6627 0 diode
R6628 N6627 N6628 10
D6628 N6628 0 diode
R6629 N6628 N6629 10
D6629 N6629 0 diode
R6630 N6629 N6630 10
D6630 N6630 0 diode
R6631 N6630 N6631 10
D6631 N6631 0 diode
R6632 N6631 N6632 10
D6632 N6632 0 diode
R6633 N6632 N6633 10
D6633 N6633 0 diode
R6634 N6633 N6634 10
D6634 N6634 0 diode
R6635 N6634 N6635 10
D6635 N6635 0 diode
R6636 N6635 N6636 10
D6636 N6636 0 diode
R6637 N6636 N6637 10
D6637 N6637 0 diode
R6638 N6637 N6638 10
D6638 N6638 0 diode
R6639 N6638 N6639 10
D6639 N6639 0 diode
R6640 N6639 N6640 10
D6640 N6640 0 diode
R6641 N6640 N6641 10
D6641 N6641 0 diode
R6642 N6641 N6642 10
D6642 N6642 0 diode
R6643 N6642 N6643 10
D6643 N6643 0 diode
R6644 N6643 N6644 10
D6644 N6644 0 diode
R6645 N6644 N6645 10
D6645 N6645 0 diode
R6646 N6645 N6646 10
D6646 N6646 0 diode
R6647 N6646 N6647 10
D6647 N6647 0 diode
R6648 N6647 N6648 10
D6648 N6648 0 diode
R6649 N6648 N6649 10
D6649 N6649 0 diode
R6650 N6649 N6650 10
D6650 N6650 0 diode
R6651 N6650 N6651 10
D6651 N6651 0 diode
R6652 N6651 N6652 10
D6652 N6652 0 diode
R6653 N6652 N6653 10
D6653 N6653 0 diode
R6654 N6653 N6654 10
D6654 N6654 0 diode
R6655 N6654 N6655 10
D6655 N6655 0 diode
R6656 N6655 N6656 10
D6656 N6656 0 diode
R6657 N6656 N6657 10
D6657 N6657 0 diode
R6658 N6657 N6658 10
D6658 N6658 0 diode
R6659 N6658 N6659 10
D6659 N6659 0 diode
R6660 N6659 N6660 10
D6660 N6660 0 diode
R6661 N6660 N6661 10
D6661 N6661 0 diode
R6662 N6661 N6662 10
D6662 N6662 0 diode
R6663 N6662 N6663 10
D6663 N6663 0 diode
R6664 N6663 N6664 10
D6664 N6664 0 diode
R6665 N6664 N6665 10
D6665 N6665 0 diode
R6666 N6665 N6666 10
D6666 N6666 0 diode
R6667 N6666 N6667 10
D6667 N6667 0 diode
R6668 N6667 N6668 10
D6668 N6668 0 diode
R6669 N6668 N6669 10
D6669 N6669 0 diode
R6670 N6669 N6670 10
D6670 N6670 0 diode
R6671 N6670 N6671 10
D6671 N6671 0 diode
R6672 N6671 N6672 10
D6672 N6672 0 diode
R6673 N6672 N6673 10
D6673 N6673 0 diode
R6674 N6673 N6674 10
D6674 N6674 0 diode
R6675 N6674 N6675 10
D6675 N6675 0 diode
R6676 N6675 N6676 10
D6676 N6676 0 diode
R6677 N6676 N6677 10
D6677 N6677 0 diode
R6678 N6677 N6678 10
D6678 N6678 0 diode
R6679 N6678 N6679 10
D6679 N6679 0 diode
R6680 N6679 N6680 10
D6680 N6680 0 diode
R6681 N6680 N6681 10
D6681 N6681 0 diode
R6682 N6681 N6682 10
D6682 N6682 0 diode
R6683 N6682 N6683 10
D6683 N6683 0 diode
R6684 N6683 N6684 10
D6684 N6684 0 diode
R6685 N6684 N6685 10
D6685 N6685 0 diode
R6686 N6685 N6686 10
D6686 N6686 0 diode
R6687 N6686 N6687 10
D6687 N6687 0 diode
R6688 N6687 N6688 10
D6688 N6688 0 diode
R6689 N6688 N6689 10
D6689 N6689 0 diode
R6690 N6689 N6690 10
D6690 N6690 0 diode
R6691 N6690 N6691 10
D6691 N6691 0 diode
R6692 N6691 N6692 10
D6692 N6692 0 diode
R6693 N6692 N6693 10
D6693 N6693 0 diode
R6694 N6693 N6694 10
D6694 N6694 0 diode
R6695 N6694 N6695 10
D6695 N6695 0 diode
R6696 N6695 N6696 10
D6696 N6696 0 diode
R6697 N6696 N6697 10
D6697 N6697 0 diode
R6698 N6697 N6698 10
D6698 N6698 0 diode
R6699 N6698 N6699 10
D6699 N6699 0 diode
R6700 N6699 N6700 10
D6700 N6700 0 diode
R6701 N6700 N6701 10
D6701 N6701 0 diode
R6702 N6701 N6702 10
D6702 N6702 0 diode
R6703 N6702 N6703 10
D6703 N6703 0 diode
R6704 N6703 N6704 10
D6704 N6704 0 diode
R6705 N6704 N6705 10
D6705 N6705 0 diode
R6706 N6705 N6706 10
D6706 N6706 0 diode
R6707 N6706 N6707 10
D6707 N6707 0 diode
R6708 N6707 N6708 10
D6708 N6708 0 diode
R6709 N6708 N6709 10
D6709 N6709 0 diode
R6710 N6709 N6710 10
D6710 N6710 0 diode
R6711 N6710 N6711 10
D6711 N6711 0 diode
R6712 N6711 N6712 10
D6712 N6712 0 diode
R6713 N6712 N6713 10
D6713 N6713 0 diode
R6714 N6713 N6714 10
D6714 N6714 0 diode
R6715 N6714 N6715 10
D6715 N6715 0 diode
R6716 N6715 N6716 10
D6716 N6716 0 diode
R6717 N6716 N6717 10
D6717 N6717 0 diode
R6718 N6717 N6718 10
D6718 N6718 0 diode
R6719 N6718 N6719 10
D6719 N6719 0 diode
R6720 N6719 N6720 10
D6720 N6720 0 diode
R6721 N6720 N6721 10
D6721 N6721 0 diode
R6722 N6721 N6722 10
D6722 N6722 0 diode
R6723 N6722 N6723 10
D6723 N6723 0 diode
R6724 N6723 N6724 10
D6724 N6724 0 diode
R6725 N6724 N6725 10
D6725 N6725 0 diode
R6726 N6725 N6726 10
D6726 N6726 0 diode
R6727 N6726 N6727 10
D6727 N6727 0 diode
R6728 N6727 N6728 10
D6728 N6728 0 diode
R6729 N6728 N6729 10
D6729 N6729 0 diode
R6730 N6729 N6730 10
D6730 N6730 0 diode
R6731 N6730 N6731 10
D6731 N6731 0 diode
R6732 N6731 N6732 10
D6732 N6732 0 diode
R6733 N6732 N6733 10
D6733 N6733 0 diode
R6734 N6733 N6734 10
D6734 N6734 0 diode
R6735 N6734 N6735 10
D6735 N6735 0 diode
R6736 N6735 N6736 10
D6736 N6736 0 diode
R6737 N6736 N6737 10
D6737 N6737 0 diode
R6738 N6737 N6738 10
D6738 N6738 0 diode
R6739 N6738 N6739 10
D6739 N6739 0 diode
R6740 N6739 N6740 10
D6740 N6740 0 diode
R6741 N6740 N6741 10
D6741 N6741 0 diode
R6742 N6741 N6742 10
D6742 N6742 0 diode
R6743 N6742 N6743 10
D6743 N6743 0 diode
R6744 N6743 N6744 10
D6744 N6744 0 diode
R6745 N6744 N6745 10
D6745 N6745 0 diode
R6746 N6745 N6746 10
D6746 N6746 0 diode
R6747 N6746 N6747 10
D6747 N6747 0 diode
R6748 N6747 N6748 10
D6748 N6748 0 diode
R6749 N6748 N6749 10
D6749 N6749 0 diode
R6750 N6749 N6750 10
D6750 N6750 0 diode
R6751 N6750 N6751 10
D6751 N6751 0 diode
R6752 N6751 N6752 10
D6752 N6752 0 diode
R6753 N6752 N6753 10
D6753 N6753 0 diode
R6754 N6753 N6754 10
D6754 N6754 0 diode
R6755 N6754 N6755 10
D6755 N6755 0 diode
R6756 N6755 N6756 10
D6756 N6756 0 diode
R6757 N6756 N6757 10
D6757 N6757 0 diode
R6758 N6757 N6758 10
D6758 N6758 0 diode
R6759 N6758 N6759 10
D6759 N6759 0 diode
R6760 N6759 N6760 10
D6760 N6760 0 diode
R6761 N6760 N6761 10
D6761 N6761 0 diode
R6762 N6761 N6762 10
D6762 N6762 0 diode
R6763 N6762 N6763 10
D6763 N6763 0 diode
R6764 N6763 N6764 10
D6764 N6764 0 diode
R6765 N6764 N6765 10
D6765 N6765 0 diode
R6766 N6765 N6766 10
D6766 N6766 0 diode
R6767 N6766 N6767 10
D6767 N6767 0 diode
R6768 N6767 N6768 10
D6768 N6768 0 diode
R6769 N6768 N6769 10
D6769 N6769 0 diode
R6770 N6769 N6770 10
D6770 N6770 0 diode
R6771 N6770 N6771 10
D6771 N6771 0 diode
R6772 N6771 N6772 10
D6772 N6772 0 diode
R6773 N6772 N6773 10
D6773 N6773 0 diode
R6774 N6773 N6774 10
D6774 N6774 0 diode
R6775 N6774 N6775 10
D6775 N6775 0 diode
R6776 N6775 N6776 10
D6776 N6776 0 diode
R6777 N6776 N6777 10
D6777 N6777 0 diode
R6778 N6777 N6778 10
D6778 N6778 0 diode
R6779 N6778 N6779 10
D6779 N6779 0 diode
R6780 N6779 N6780 10
D6780 N6780 0 diode
R6781 N6780 N6781 10
D6781 N6781 0 diode
R6782 N6781 N6782 10
D6782 N6782 0 diode
R6783 N6782 N6783 10
D6783 N6783 0 diode
R6784 N6783 N6784 10
D6784 N6784 0 diode
R6785 N6784 N6785 10
D6785 N6785 0 diode
R6786 N6785 N6786 10
D6786 N6786 0 diode
R6787 N6786 N6787 10
D6787 N6787 0 diode
R6788 N6787 N6788 10
D6788 N6788 0 diode
R6789 N6788 N6789 10
D6789 N6789 0 diode
R6790 N6789 N6790 10
D6790 N6790 0 diode
R6791 N6790 N6791 10
D6791 N6791 0 diode
R6792 N6791 N6792 10
D6792 N6792 0 diode
R6793 N6792 N6793 10
D6793 N6793 0 diode
R6794 N6793 N6794 10
D6794 N6794 0 diode
R6795 N6794 N6795 10
D6795 N6795 0 diode
R6796 N6795 N6796 10
D6796 N6796 0 diode
R6797 N6796 N6797 10
D6797 N6797 0 diode
R6798 N6797 N6798 10
D6798 N6798 0 diode
R6799 N6798 N6799 10
D6799 N6799 0 diode
R6800 N6799 N6800 10
D6800 N6800 0 diode
R6801 N6800 N6801 10
D6801 N6801 0 diode
R6802 N6801 N6802 10
D6802 N6802 0 diode
R6803 N6802 N6803 10
D6803 N6803 0 diode
R6804 N6803 N6804 10
D6804 N6804 0 diode
R6805 N6804 N6805 10
D6805 N6805 0 diode
R6806 N6805 N6806 10
D6806 N6806 0 diode
R6807 N6806 N6807 10
D6807 N6807 0 diode
R6808 N6807 N6808 10
D6808 N6808 0 diode
R6809 N6808 N6809 10
D6809 N6809 0 diode
R6810 N6809 N6810 10
D6810 N6810 0 diode
R6811 N6810 N6811 10
D6811 N6811 0 diode
R6812 N6811 N6812 10
D6812 N6812 0 diode
R6813 N6812 N6813 10
D6813 N6813 0 diode
R6814 N6813 N6814 10
D6814 N6814 0 diode
R6815 N6814 N6815 10
D6815 N6815 0 diode
R6816 N6815 N6816 10
D6816 N6816 0 diode
R6817 N6816 N6817 10
D6817 N6817 0 diode
R6818 N6817 N6818 10
D6818 N6818 0 diode
R6819 N6818 N6819 10
D6819 N6819 0 diode
R6820 N6819 N6820 10
D6820 N6820 0 diode
R6821 N6820 N6821 10
D6821 N6821 0 diode
R6822 N6821 N6822 10
D6822 N6822 0 diode
R6823 N6822 N6823 10
D6823 N6823 0 diode
R6824 N6823 N6824 10
D6824 N6824 0 diode
R6825 N6824 N6825 10
D6825 N6825 0 diode
R6826 N6825 N6826 10
D6826 N6826 0 diode
R6827 N6826 N6827 10
D6827 N6827 0 diode
R6828 N6827 N6828 10
D6828 N6828 0 diode
R6829 N6828 N6829 10
D6829 N6829 0 diode
R6830 N6829 N6830 10
D6830 N6830 0 diode
R6831 N6830 N6831 10
D6831 N6831 0 diode
R6832 N6831 N6832 10
D6832 N6832 0 diode
R6833 N6832 N6833 10
D6833 N6833 0 diode
R6834 N6833 N6834 10
D6834 N6834 0 diode
R6835 N6834 N6835 10
D6835 N6835 0 diode
R6836 N6835 N6836 10
D6836 N6836 0 diode
R6837 N6836 N6837 10
D6837 N6837 0 diode
R6838 N6837 N6838 10
D6838 N6838 0 diode
R6839 N6838 N6839 10
D6839 N6839 0 diode
R6840 N6839 N6840 10
D6840 N6840 0 diode
R6841 N6840 N6841 10
D6841 N6841 0 diode
R6842 N6841 N6842 10
D6842 N6842 0 diode
R6843 N6842 N6843 10
D6843 N6843 0 diode
R6844 N6843 N6844 10
D6844 N6844 0 diode
R6845 N6844 N6845 10
D6845 N6845 0 diode
R6846 N6845 N6846 10
D6846 N6846 0 diode
R6847 N6846 N6847 10
D6847 N6847 0 diode
R6848 N6847 N6848 10
D6848 N6848 0 diode
R6849 N6848 N6849 10
D6849 N6849 0 diode
R6850 N6849 N6850 10
D6850 N6850 0 diode
R6851 N6850 N6851 10
D6851 N6851 0 diode
R6852 N6851 N6852 10
D6852 N6852 0 diode
R6853 N6852 N6853 10
D6853 N6853 0 diode
R6854 N6853 N6854 10
D6854 N6854 0 diode
R6855 N6854 N6855 10
D6855 N6855 0 diode
R6856 N6855 N6856 10
D6856 N6856 0 diode
R6857 N6856 N6857 10
D6857 N6857 0 diode
R6858 N6857 N6858 10
D6858 N6858 0 diode
R6859 N6858 N6859 10
D6859 N6859 0 diode
R6860 N6859 N6860 10
D6860 N6860 0 diode
R6861 N6860 N6861 10
D6861 N6861 0 diode
R6862 N6861 N6862 10
D6862 N6862 0 diode
R6863 N6862 N6863 10
D6863 N6863 0 diode
R6864 N6863 N6864 10
D6864 N6864 0 diode
R6865 N6864 N6865 10
D6865 N6865 0 diode
R6866 N6865 N6866 10
D6866 N6866 0 diode
R6867 N6866 N6867 10
D6867 N6867 0 diode
R6868 N6867 N6868 10
D6868 N6868 0 diode
R6869 N6868 N6869 10
D6869 N6869 0 diode
R6870 N6869 N6870 10
D6870 N6870 0 diode
R6871 N6870 N6871 10
D6871 N6871 0 diode
R6872 N6871 N6872 10
D6872 N6872 0 diode
R6873 N6872 N6873 10
D6873 N6873 0 diode
R6874 N6873 N6874 10
D6874 N6874 0 diode
R6875 N6874 N6875 10
D6875 N6875 0 diode
R6876 N6875 N6876 10
D6876 N6876 0 diode
R6877 N6876 N6877 10
D6877 N6877 0 diode
R6878 N6877 N6878 10
D6878 N6878 0 diode
R6879 N6878 N6879 10
D6879 N6879 0 diode
R6880 N6879 N6880 10
D6880 N6880 0 diode
R6881 N6880 N6881 10
D6881 N6881 0 diode
R6882 N6881 N6882 10
D6882 N6882 0 diode
R6883 N6882 N6883 10
D6883 N6883 0 diode
R6884 N6883 N6884 10
D6884 N6884 0 diode
R6885 N6884 N6885 10
D6885 N6885 0 diode
R6886 N6885 N6886 10
D6886 N6886 0 diode
R6887 N6886 N6887 10
D6887 N6887 0 diode
R6888 N6887 N6888 10
D6888 N6888 0 diode
R6889 N6888 N6889 10
D6889 N6889 0 diode
R6890 N6889 N6890 10
D6890 N6890 0 diode
R6891 N6890 N6891 10
D6891 N6891 0 diode
R6892 N6891 N6892 10
D6892 N6892 0 diode
R6893 N6892 N6893 10
D6893 N6893 0 diode
R6894 N6893 N6894 10
D6894 N6894 0 diode
R6895 N6894 N6895 10
D6895 N6895 0 diode
R6896 N6895 N6896 10
D6896 N6896 0 diode
R6897 N6896 N6897 10
D6897 N6897 0 diode
R6898 N6897 N6898 10
D6898 N6898 0 diode
R6899 N6898 N6899 10
D6899 N6899 0 diode
R6900 N6899 N6900 10
D6900 N6900 0 diode
R6901 N6900 N6901 10
D6901 N6901 0 diode
R6902 N6901 N6902 10
D6902 N6902 0 diode
R6903 N6902 N6903 10
D6903 N6903 0 diode
R6904 N6903 N6904 10
D6904 N6904 0 diode
R6905 N6904 N6905 10
D6905 N6905 0 diode
R6906 N6905 N6906 10
D6906 N6906 0 diode
R6907 N6906 N6907 10
D6907 N6907 0 diode
R6908 N6907 N6908 10
D6908 N6908 0 diode
R6909 N6908 N6909 10
D6909 N6909 0 diode
R6910 N6909 N6910 10
D6910 N6910 0 diode
R6911 N6910 N6911 10
D6911 N6911 0 diode
R6912 N6911 N6912 10
D6912 N6912 0 diode
R6913 N6912 N6913 10
D6913 N6913 0 diode
R6914 N6913 N6914 10
D6914 N6914 0 diode
R6915 N6914 N6915 10
D6915 N6915 0 diode
R6916 N6915 N6916 10
D6916 N6916 0 diode
R6917 N6916 N6917 10
D6917 N6917 0 diode
R6918 N6917 N6918 10
D6918 N6918 0 diode
R6919 N6918 N6919 10
D6919 N6919 0 diode
R6920 N6919 N6920 10
D6920 N6920 0 diode
R6921 N6920 N6921 10
D6921 N6921 0 diode
R6922 N6921 N6922 10
D6922 N6922 0 diode
R6923 N6922 N6923 10
D6923 N6923 0 diode
R6924 N6923 N6924 10
D6924 N6924 0 diode
R6925 N6924 N6925 10
D6925 N6925 0 diode
R6926 N6925 N6926 10
D6926 N6926 0 diode
R6927 N6926 N6927 10
D6927 N6927 0 diode
R6928 N6927 N6928 10
D6928 N6928 0 diode
R6929 N6928 N6929 10
D6929 N6929 0 diode
R6930 N6929 N6930 10
D6930 N6930 0 diode
R6931 N6930 N6931 10
D6931 N6931 0 diode
R6932 N6931 N6932 10
D6932 N6932 0 diode
R6933 N6932 N6933 10
D6933 N6933 0 diode
R6934 N6933 N6934 10
D6934 N6934 0 diode
R6935 N6934 N6935 10
D6935 N6935 0 diode
R6936 N6935 N6936 10
D6936 N6936 0 diode
R6937 N6936 N6937 10
D6937 N6937 0 diode
R6938 N6937 N6938 10
D6938 N6938 0 diode
R6939 N6938 N6939 10
D6939 N6939 0 diode
R6940 N6939 N6940 10
D6940 N6940 0 diode
R6941 N6940 N6941 10
D6941 N6941 0 diode
R6942 N6941 N6942 10
D6942 N6942 0 diode
R6943 N6942 N6943 10
D6943 N6943 0 diode
R6944 N6943 N6944 10
D6944 N6944 0 diode
R6945 N6944 N6945 10
D6945 N6945 0 diode
R6946 N6945 N6946 10
D6946 N6946 0 diode
R6947 N6946 N6947 10
D6947 N6947 0 diode
R6948 N6947 N6948 10
D6948 N6948 0 diode
R6949 N6948 N6949 10
D6949 N6949 0 diode
R6950 N6949 N6950 10
D6950 N6950 0 diode
R6951 N6950 N6951 10
D6951 N6951 0 diode
R6952 N6951 N6952 10
D6952 N6952 0 diode
R6953 N6952 N6953 10
D6953 N6953 0 diode
R6954 N6953 N6954 10
D6954 N6954 0 diode
R6955 N6954 N6955 10
D6955 N6955 0 diode
R6956 N6955 N6956 10
D6956 N6956 0 diode
R6957 N6956 N6957 10
D6957 N6957 0 diode
R6958 N6957 N6958 10
D6958 N6958 0 diode
R6959 N6958 N6959 10
D6959 N6959 0 diode
R6960 N6959 N6960 10
D6960 N6960 0 diode
R6961 N6960 N6961 10
D6961 N6961 0 diode
R6962 N6961 N6962 10
D6962 N6962 0 diode
R6963 N6962 N6963 10
D6963 N6963 0 diode
R6964 N6963 N6964 10
D6964 N6964 0 diode
R6965 N6964 N6965 10
D6965 N6965 0 diode
R6966 N6965 N6966 10
D6966 N6966 0 diode
R6967 N6966 N6967 10
D6967 N6967 0 diode
R6968 N6967 N6968 10
D6968 N6968 0 diode
R6969 N6968 N6969 10
D6969 N6969 0 diode
R6970 N6969 N6970 10
D6970 N6970 0 diode
R6971 N6970 N6971 10
D6971 N6971 0 diode
R6972 N6971 N6972 10
D6972 N6972 0 diode
R6973 N6972 N6973 10
D6973 N6973 0 diode
R6974 N6973 N6974 10
D6974 N6974 0 diode
R6975 N6974 N6975 10
D6975 N6975 0 diode
R6976 N6975 N6976 10
D6976 N6976 0 diode
R6977 N6976 N6977 10
D6977 N6977 0 diode
R6978 N6977 N6978 10
D6978 N6978 0 diode
R6979 N6978 N6979 10
D6979 N6979 0 diode
R6980 N6979 N6980 10
D6980 N6980 0 diode
R6981 N6980 N6981 10
D6981 N6981 0 diode
R6982 N6981 N6982 10
D6982 N6982 0 diode
R6983 N6982 N6983 10
D6983 N6983 0 diode
R6984 N6983 N6984 10
D6984 N6984 0 diode
R6985 N6984 N6985 10
D6985 N6985 0 diode
R6986 N6985 N6986 10
D6986 N6986 0 diode
R6987 N6986 N6987 10
D6987 N6987 0 diode
R6988 N6987 N6988 10
D6988 N6988 0 diode
R6989 N6988 N6989 10
D6989 N6989 0 diode
R6990 N6989 N6990 10
D6990 N6990 0 diode
R6991 N6990 N6991 10
D6991 N6991 0 diode
R6992 N6991 N6992 10
D6992 N6992 0 diode
R6993 N6992 N6993 10
D6993 N6993 0 diode
R6994 N6993 N6994 10
D6994 N6994 0 diode
R6995 N6994 N6995 10
D6995 N6995 0 diode
R6996 N6995 N6996 10
D6996 N6996 0 diode
R6997 N6996 N6997 10
D6997 N6997 0 diode
R6998 N6997 N6998 10
D6998 N6998 0 diode
R6999 N6998 N6999 10
D6999 N6999 0 diode
R7000 N6999 N7000 10
D7000 N7000 0 diode
R7001 N7000 N7001 10
D7001 N7001 0 diode
R7002 N7001 N7002 10
D7002 N7002 0 diode
R7003 N7002 N7003 10
D7003 N7003 0 diode
R7004 N7003 N7004 10
D7004 N7004 0 diode
R7005 N7004 N7005 10
D7005 N7005 0 diode
R7006 N7005 N7006 10
D7006 N7006 0 diode
R7007 N7006 N7007 10
D7007 N7007 0 diode
R7008 N7007 N7008 10
D7008 N7008 0 diode
R7009 N7008 N7009 10
D7009 N7009 0 diode
R7010 N7009 N7010 10
D7010 N7010 0 diode
R7011 N7010 N7011 10
D7011 N7011 0 diode
R7012 N7011 N7012 10
D7012 N7012 0 diode
R7013 N7012 N7013 10
D7013 N7013 0 diode
R7014 N7013 N7014 10
D7014 N7014 0 diode
R7015 N7014 N7015 10
D7015 N7015 0 diode
R7016 N7015 N7016 10
D7016 N7016 0 diode
R7017 N7016 N7017 10
D7017 N7017 0 diode
R7018 N7017 N7018 10
D7018 N7018 0 diode
R7019 N7018 N7019 10
D7019 N7019 0 diode
R7020 N7019 N7020 10
D7020 N7020 0 diode
R7021 N7020 N7021 10
D7021 N7021 0 diode
R7022 N7021 N7022 10
D7022 N7022 0 diode
R7023 N7022 N7023 10
D7023 N7023 0 diode
R7024 N7023 N7024 10
D7024 N7024 0 diode
R7025 N7024 N7025 10
D7025 N7025 0 diode
R7026 N7025 N7026 10
D7026 N7026 0 diode
R7027 N7026 N7027 10
D7027 N7027 0 diode
R7028 N7027 N7028 10
D7028 N7028 0 diode
R7029 N7028 N7029 10
D7029 N7029 0 diode
R7030 N7029 N7030 10
D7030 N7030 0 diode
R7031 N7030 N7031 10
D7031 N7031 0 diode
R7032 N7031 N7032 10
D7032 N7032 0 diode
R7033 N7032 N7033 10
D7033 N7033 0 diode
R7034 N7033 N7034 10
D7034 N7034 0 diode
R7035 N7034 N7035 10
D7035 N7035 0 diode
R7036 N7035 N7036 10
D7036 N7036 0 diode
R7037 N7036 N7037 10
D7037 N7037 0 diode
R7038 N7037 N7038 10
D7038 N7038 0 diode
R7039 N7038 N7039 10
D7039 N7039 0 diode
R7040 N7039 N7040 10
D7040 N7040 0 diode
R7041 N7040 N7041 10
D7041 N7041 0 diode
R7042 N7041 N7042 10
D7042 N7042 0 diode
R7043 N7042 N7043 10
D7043 N7043 0 diode
R7044 N7043 N7044 10
D7044 N7044 0 diode
R7045 N7044 N7045 10
D7045 N7045 0 diode
R7046 N7045 N7046 10
D7046 N7046 0 diode
R7047 N7046 N7047 10
D7047 N7047 0 diode
R7048 N7047 N7048 10
D7048 N7048 0 diode
R7049 N7048 N7049 10
D7049 N7049 0 diode
R7050 N7049 N7050 10
D7050 N7050 0 diode
R7051 N7050 N7051 10
D7051 N7051 0 diode
R7052 N7051 N7052 10
D7052 N7052 0 diode
R7053 N7052 N7053 10
D7053 N7053 0 diode
R7054 N7053 N7054 10
D7054 N7054 0 diode
R7055 N7054 N7055 10
D7055 N7055 0 diode
R7056 N7055 N7056 10
D7056 N7056 0 diode
R7057 N7056 N7057 10
D7057 N7057 0 diode
R7058 N7057 N7058 10
D7058 N7058 0 diode
R7059 N7058 N7059 10
D7059 N7059 0 diode
R7060 N7059 N7060 10
D7060 N7060 0 diode
R7061 N7060 N7061 10
D7061 N7061 0 diode
R7062 N7061 N7062 10
D7062 N7062 0 diode
R7063 N7062 N7063 10
D7063 N7063 0 diode
R7064 N7063 N7064 10
D7064 N7064 0 diode
R7065 N7064 N7065 10
D7065 N7065 0 diode
R7066 N7065 N7066 10
D7066 N7066 0 diode
R7067 N7066 N7067 10
D7067 N7067 0 diode
R7068 N7067 N7068 10
D7068 N7068 0 diode
R7069 N7068 N7069 10
D7069 N7069 0 diode
R7070 N7069 N7070 10
D7070 N7070 0 diode
R7071 N7070 N7071 10
D7071 N7071 0 diode
R7072 N7071 N7072 10
D7072 N7072 0 diode
R7073 N7072 N7073 10
D7073 N7073 0 diode
R7074 N7073 N7074 10
D7074 N7074 0 diode
R7075 N7074 N7075 10
D7075 N7075 0 diode
R7076 N7075 N7076 10
D7076 N7076 0 diode
R7077 N7076 N7077 10
D7077 N7077 0 diode
R7078 N7077 N7078 10
D7078 N7078 0 diode
R7079 N7078 N7079 10
D7079 N7079 0 diode
R7080 N7079 N7080 10
D7080 N7080 0 diode
R7081 N7080 N7081 10
D7081 N7081 0 diode
R7082 N7081 N7082 10
D7082 N7082 0 diode
R7083 N7082 N7083 10
D7083 N7083 0 diode
R7084 N7083 N7084 10
D7084 N7084 0 diode
R7085 N7084 N7085 10
D7085 N7085 0 diode
R7086 N7085 N7086 10
D7086 N7086 0 diode
R7087 N7086 N7087 10
D7087 N7087 0 diode
R7088 N7087 N7088 10
D7088 N7088 0 diode
R7089 N7088 N7089 10
D7089 N7089 0 diode
R7090 N7089 N7090 10
D7090 N7090 0 diode
R7091 N7090 N7091 10
D7091 N7091 0 diode
R7092 N7091 N7092 10
D7092 N7092 0 diode
R7093 N7092 N7093 10
D7093 N7093 0 diode
R7094 N7093 N7094 10
D7094 N7094 0 diode
R7095 N7094 N7095 10
D7095 N7095 0 diode
R7096 N7095 N7096 10
D7096 N7096 0 diode
R7097 N7096 N7097 10
D7097 N7097 0 diode
R7098 N7097 N7098 10
D7098 N7098 0 diode
R7099 N7098 N7099 10
D7099 N7099 0 diode
R7100 N7099 N7100 10
D7100 N7100 0 diode
R7101 N7100 N7101 10
D7101 N7101 0 diode
R7102 N7101 N7102 10
D7102 N7102 0 diode
R7103 N7102 N7103 10
D7103 N7103 0 diode
R7104 N7103 N7104 10
D7104 N7104 0 diode
R7105 N7104 N7105 10
D7105 N7105 0 diode
R7106 N7105 N7106 10
D7106 N7106 0 diode
R7107 N7106 N7107 10
D7107 N7107 0 diode
R7108 N7107 N7108 10
D7108 N7108 0 diode
R7109 N7108 N7109 10
D7109 N7109 0 diode
R7110 N7109 N7110 10
D7110 N7110 0 diode
R7111 N7110 N7111 10
D7111 N7111 0 diode
R7112 N7111 N7112 10
D7112 N7112 0 diode
R7113 N7112 N7113 10
D7113 N7113 0 diode
R7114 N7113 N7114 10
D7114 N7114 0 diode
R7115 N7114 N7115 10
D7115 N7115 0 diode
R7116 N7115 N7116 10
D7116 N7116 0 diode
R7117 N7116 N7117 10
D7117 N7117 0 diode
R7118 N7117 N7118 10
D7118 N7118 0 diode
R7119 N7118 N7119 10
D7119 N7119 0 diode
R7120 N7119 N7120 10
D7120 N7120 0 diode
R7121 N7120 N7121 10
D7121 N7121 0 diode
R7122 N7121 N7122 10
D7122 N7122 0 diode
R7123 N7122 N7123 10
D7123 N7123 0 diode
R7124 N7123 N7124 10
D7124 N7124 0 diode
R7125 N7124 N7125 10
D7125 N7125 0 diode
R7126 N7125 N7126 10
D7126 N7126 0 diode
R7127 N7126 N7127 10
D7127 N7127 0 diode
R7128 N7127 N7128 10
D7128 N7128 0 diode
R7129 N7128 N7129 10
D7129 N7129 0 diode
R7130 N7129 N7130 10
D7130 N7130 0 diode
R7131 N7130 N7131 10
D7131 N7131 0 diode
R7132 N7131 N7132 10
D7132 N7132 0 diode
R7133 N7132 N7133 10
D7133 N7133 0 diode
R7134 N7133 N7134 10
D7134 N7134 0 diode
R7135 N7134 N7135 10
D7135 N7135 0 diode
R7136 N7135 N7136 10
D7136 N7136 0 diode
R7137 N7136 N7137 10
D7137 N7137 0 diode
R7138 N7137 N7138 10
D7138 N7138 0 diode
R7139 N7138 N7139 10
D7139 N7139 0 diode
R7140 N7139 N7140 10
D7140 N7140 0 diode
R7141 N7140 N7141 10
D7141 N7141 0 diode
R7142 N7141 N7142 10
D7142 N7142 0 diode
R7143 N7142 N7143 10
D7143 N7143 0 diode
R7144 N7143 N7144 10
D7144 N7144 0 diode
R7145 N7144 N7145 10
D7145 N7145 0 diode
R7146 N7145 N7146 10
D7146 N7146 0 diode
R7147 N7146 N7147 10
D7147 N7147 0 diode
R7148 N7147 N7148 10
D7148 N7148 0 diode
R7149 N7148 N7149 10
D7149 N7149 0 diode
R7150 N7149 N7150 10
D7150 N7150 0 diode
R7151 N7150 N7151 10
D7151 N7151 0 diode
R7152 N7151 N7152 10
D7152 N7152 0 diode
R7153 N7152 N7153 10
D7153 N7153 0 diode
R7154 N7153 N7154 10
D7154 N7154 0 diode
R7155 N7154 N7155 10
D7155 N7155 0 diode
R7156 N7155 N7156 10
D7156 N7156 0 diode
R7157 N7156 N7157 10
D7157 N7157 0 diode
R7158 N7157 N7158 10
D7158 N7158 0 diode
R7159 N7158 N7159 10
D7159 N7159 0 diode
R7160 N7159 N7160 10
D7160 N7160 0 diode
R7161 N7160 N7161 10
D7161 N7161 0 diode
R7162 N7161 N7162 10
D7162 N7162 0 diode
R7163 N7162 N7163 10
D7163 N7163 0 diode
R7164 N7163 N7164 10
D7164 N7164 0 diode
R7165 N7164 N7165 10
D7165 N7165 0 diode
R7166 N7165 N7166 10
D7166 N7166 0 diode
R7167 N7166 N7167 10
D7167 N7167 0 diode
R7168 N7167 N7168 10
D7168 N7168 0 diode
R7169 N7168 N7169 10
D7169 N7169 0 diode
R7170 N7169 N7170 10
D7170 N7170 0 diode
R7171 N7170 N7171 10
D7171 N7171 0 diode
R7172 N7171 N7172 10
D7172 N7172 0 diode
R7173 N7172 N7173 10
D7173 N7173 0 diode
R7174 N7173 N7174 10
D7174 N7174 0 diode
R7175 N7174 N7175 10
D7175 N7175 0 diode
R7176 N7175 N7176 10
D7176 N7176 0 diode
R7177 N7176 N7177 10
D7177 N7177 0 diode
R7178 N7177 N7178 10
D7178 N7178 0 diode
R7179 N7178 N7179 10
D7179 N7179 0 diode
R7180 N7179 N7180 10
D7180 N7180 0 diode
R7181 N7180 N7181 10
D7181 N7181 0 diode
R7182 N7181 N7182 10
D7182 N7182 0 diode
R7183 N7182 N7183 10
D7183 N7183 0 diode
R7184 N7183 N7184 10
D7184 N7184 0 diode
R7185 N7184 N7185 10
D7185 N7185 0 diode
R7186 N7185 N7186 10
D7186 N7186 0 diode
R7187 N7186 N7187 10
D7187 N7187 0 diode
R7188 N7187 N7188 10
D7188 N7188 0 diode
R7189 N7188 N7189 10
D7189 N7189 0 diode
R7190 N7189 N7190 10
D7190 N7190 0 diode
R7191 N7190 N7191 10
D7191 N7191 0 diode
R7192 N7191 N7192 10
D7192 N7192 0 diode
R7193 N7192 N7193 10
D7193 N7193 0 diode
R7194 N7193 N7194 10
D7194 N7194 0 diode
R7195 N7194 N7195 10
D7195 N7195 0 diode
R7196 N7195 N7196 10
D7196 N7196 0 diode
R7197 N7196 N7197 10
D7197 N7197 0 diode
R7198 N7197 N7198 10
D7198 N7198 0 diode
R7199 N7198 N7199 10
D7199 N7199 0 diode
R7200 N7199 N7200 10
D7200 N7200 0 diode
R7201 N7200 N7201 10
D7201 N7201 0 diode
R7202 N7201 N7202 10
D7202 N7202 0 diode
R7203 N7202 N7203 10
D7203 N7203 0 diode
R7204 N7203 N7204 10
D7204 N7204 0 diode
R7205 N7204 N7205 10
D7205 N7205 0 diode
R7206 N7205 N7206 10
D7206 N7206 0 diode
R7207 N7206 N7207 10
D7207 N7207 0 diode
R7208 N7207 N7208 10
D7208 N7208 0 diode
R7209 N7208 N7209 10
D7209 N7209 0 diode
R7210 N7209 N7210 10
D7210 N7210 0 diode
R7211 N7210 N7211 10
D7211 N7211 0 diode
R7212 N7211 N7212 10
D7212 N7212 0 diode
R7213 N7212 N7213 10
D7213 N7213 0 diode
R7214 N7213 N7214 10
D7214 N7214 0 diode
R7215 N7214 N7215 10
D7215 N7215 0 diode
R7216 N7215 N7216 10
D7216 N7216 0 diode
R7217 N7216 N7217 10
D7217 N7217 0 diode
R7218 N7217 N7218 10
D7218 N7218 0 diode
R7219 N7218 N7219 10
D7219 N7219 0 diode
R7220 N7219 N7220 10
D7220 N7220 0 diode
R7221 N7220 N7221 10
D7221 N7221 0 diode
R7222 N7221 N7222 10
D7222 N7222 0 diode
R7223 N7222 N7223 10
D7223 N7223 0 diode
R7224 N7223 N7224 10
D7224 N7224 0 diode
R7225 N7224 N7225 10
D7225 N7225 0 diode
R7226 N7225 N7226 10
D7226 N7226 0 diode
R7227 N7226 N7227 10
D7227 N7227 0 diode
R7228 N7227 N7228 10
D7228 N7228 0 diode
R7229 N7228 N7229 10
D7229 N7229 0 diode
R7230 N7229 N7230 10
D7230 N7230 0 diode
R7231 N7230 N7231 10
D7231 N7231 0 diode
R7232 N7231 N7232 10
D7232 N7232 0 diode
R7233 N7232 N7233 10
D7233 N7233 0 diode
R7234 N7233 N7234 10
D7234 N7234 0 diode
R7235 N7234 N7235 10
D7235 N7235 0 diode
R7236 N7235 N7236 10
D7236 N7236 0 diode
R7237 N7236 N7237 10
D7237 N7237 0 diode
R7238 N7237 N7238 10
D7238 N7238 0 diode
R7239 N7238 N7239 10
D7239 N7239 0 diode
R7240 N7239 N7240 10
D7240 N7240 0 diode
R7241 N7240 N7241 10
D7241 N7241 0 diode
R7242 N7241 N7242 10
D7242 N7242 0 diode
R7243 N7242 N7243 10
D7243 N7243 0 diode
R7244 N7243 N7244 10
D7244 N7244 0 diode
R7245 N7244 N7245 10
D7245 N7245 0 diode
R7246 N7245 N7246 10
D7246 N7246 0 diode
R7247 N7246 N7247 10
D7247 N7247 0 diode
R7248 N7247 N7248 10
D7248 N7248 0 diode
R7249 N7248 N7249 10
D7249 N7249 0 diode
R7250 N7249 N7250 10
D7250 N7250 0 diode
R7251 N7250 N7251 10
D7251 N7251 0 diode
R7252 N7251 N7252 10
D7252 N7252 0 diode
R7253 N7252 N7253 10
D7253 N7253 0 diode
R7254 N7253 N7254 10
D7254 N7254 0 diode
R7255 N7254 N7255 10
D7255 N7255 0 diode
R7256 N7255 N7256 10
D7256 N7256 0 diode
R7257 N7256 N7257 10
D7257 N7257 0 diode
R7258 N7257 N7258 10
D7258 N7258 0 diode
R7259 N7258 N7259 10
D7259 N7259 0 diode
R7260 N7259 N7260 10
D7260 N7260 0 diode
R7261 N7260 N7261 10
D7261 N7261 0 diode
R7262 N7261 N7262 10
D7262 N7262 0 diode
R7263 N7262 N7263 10
D7263 N7263 0 diode
R7264 N7263 N7264 10
D7264 N7264 0 diode
R7265 N7264 N7265 10
D7265 N7265 0 diode
R7266 N7265 N7266 10
D7266 N7266 0 diode
R7267 N7266 N7267 10
D7267 N7267 0 diode
R7268 N7267 N7268 10
D7268 N7268 0 diode
R7269 N7268 N7269 10
D7269 N7269 0 diode
R7270 N7269 N7270 10
D7270 N7270 0 diode
R7271 N7270 N7271 10
D7271 N7271 0 diode
R7272 N7271 N7272 10
D7272 N7272 0 diode
R7273 N7272 N7273 10
D7273 N7273 0 diode
R7274 N7273 N7274 10
D7274 N7274 0 diode
R7275 N7274 N7275 10
D7275 N7275 0 diode
R7276 N7275 N7276 10
D7276 N7276 0 diode
R7277 N7276 N7277 10
D7277 N7277 0 diode
R7278 N7277 N7278 10
D7278 N7278 0 diode
R7279 N7278 N7279 10
D7279 N7279 0 diode
R7280 N7279 N7280 10
D7280 N7280 0 diode
R7281 N7280 N7281 10
D7281 N7281 0 diode
R7282 N7281 N7282 10
D7282 N7282 0 diode
R7283 N7282 N7283 10
D7283 N7283 0 diode
R7284 N7283 N7284 10
D7284 N7284 0 diode
R7285 N7284 N7285 10
D7285 N7285 0 diode
R7286 N7285 N7286 10
D7286 N7286 0 diode
R7287 N7286 N7287 10
D7287 N7287 0 diode
R7288 N7287 N7288 10
D7288 N7288 0 diode
R7289 N7288 N7289 10
D7289 N7289 0 diode
R7290 N7289 N7290 10
D7290 N7290 0 diode
R7291 N7290 N7291 10
D7291 N7291 0 diode
R7292 N7291 N7292 10
D7292 N7292 0 diode
R7293 N7292 N7293 10
D7293 N7293 0 diode
R7294 N7293 N7294 10
D7294 N7294 0 diode
R7295 N7294 N7295 10
D7295 N7295 0 diode
R7296 N7295 N7296 10
D7296 N7296 0 diode
R7297 N7296 N7297 10
D7297 N7297 0 diode
R7298 N7297 N7298 10
D7298 N7298 0 diode
R7299 N7298 N7299 10
D7299 N7299 0 diode
R7300 N7299 N7300 10
D7300 N7300 0 diode
R7301 N7300 N7301 10
D7301 N7301 0 diode
R7302 N7301 N7302 10
D7302 N7302 0 diode
R7303 N7302 N7303 10
D7303 N7303 0 diode
R7304 N7303 N7304 10
D7304 N7304 0 diode
R7305 N7304 N7305 10
D7305 N7305 0 diode
R7306 N7305 N7306 10
D7306 N7306 0 diode
R7307 N7306 N7307 10
D7307 N7307 0 diode
R7308 N7307 N7308 10
D7308 N7308 0 diode
R7309 N7308 N7309 10
D7309 N7309 0 diode
R7310 N7309 N7310 10
D7310 N7310 0 diode
R7311 N7310 N7311 10
D7311 N7311 0 diode
R7312 N7311 N7312 10
D7312 N7312 0 diode
R7313 N7312 N7313 10
D7313 N7313 0 diode
R7314 N7313 N7314 10
D7314 N7314 0 diode
R7315 N7314 N7315 10
D7315 N7315 0 diode
R7316 N7315 N7316 10
D7316 N7316 0 diode
R7317 N7316 N7317 10
D7317 N7317 0 diode
R7318 N7317 N7318 10
D7318 N7318 0 diode
R7319 N7318 N7319 10
D7319 N7319 0 diode
R7320 N7319 N7320 10
D7320 N7320 0 diode
R7321 N7320 N7321 10
D7321 N7321 0 diode
R7322 N7321 N7322 10
D7322 N7322 0 diode
R7323 N7322 N7323 10
D7323 N7323 0 diode
R7324 N7323 N7324 10
D7324 N7324 0 diode
R7325 N7324 N7325 10
D7325 N7325 0 diode
R7326 N7325 N7326 10
D7326 N7326 0 diode
R7327 N7326 N7327 10
D7327 N7327 0 diode
R7328 N7327 N7328 10
D7328 N7328 0 diode
R7329 N7328 N7329 10
D7329 N7329 0 diode
R7330 N7329 N7330 10
D7330 N7330 0 diode
R7331 N7330 N7331 10
D7331 N7331 0 diode
R7332 N7331 N7332 10
D7332 N7332 0 diode
R7333 N7332 N7333 10
D7333 N7333 0 diode
R7334 N7333 N7334 10
D7334 N7334 0 diode
R7335 N7334 N7335 10
D7335 N7335 0 diode
R7336 N7335 N7336 10
D7336 N7336 0 diode
R7337 N7336 N7337 10
D7337 N7337 0 diode
R7338 N7337 N7338 10
D7338 N7338 0 diode
R7339 N7338 N7339 10
D7339 N7339 0 diode
R7340 N7339 N7340 10
D7340 N7340 0 diode
R7341 N7340 N7341 10
D7341 N7341 0 diode
R7342 N7341 N7342 10
D7342 N7342 0 diode
R7343 N7342 N7343 10
D7343 N7343 0 diode
R7344 N7343 N7344 10
D7344 N7344 0 diode
R7345 N7344 N7345 10
D7345 N7345 0 diode
R7346 N7345 N7346 10
D7346 N7346 0 diode
R7347 N7346 N7347 10
D7347 N7347 0 diode
R7348 N7347 N7348 10
D7348 N7348 0 diode
R7349 N7348 N7349 10
D7349 N7349 0 diode
R7350 N7349 N7350 10
D7350 N7350 0 diode
R7351 N7350 N7351 10
D7351 N7351 0 diode
R7352 N7351 N7352 10
D7352 N7352 0 diode
R7353 N7352 N7353 10
D7353 N7353 0 diode
R7354 N7353 N7354 10
D7354 N7354 0 diode
R7355 N7354 N7355 10
D7355 N7355 0 diode
R7356 N7355 N7356 10
D7356 N7356 0 diode
R7357 N7356 N7357 10
D7357 N7357 0 diode
R7358 N7357 N7358 10
D7358 N7358 0 diode
R7359 N7358 N7359 10
D7359 N7359 0 diode
R7360 N7359 N7360 10
D7360 N7360 0 diode
R7361 N7360 N7361 10
D7361 N7361 0 diode
R7362 N7361 N7362 10
D7362 N7362 0 diode
R7363 N7362 N7363 10
D7363 N7363 0 diode
R7364 N7363 N7364 10
D7364 N7364 0 diode
R7365 N7364 N7365 10
D7365 N7365 0 diode
R7366 N7365 N7366 10
D7366 N7366 0 diode
R7367 N7366 N7367 10
D7367 N7367 0 diode
R7368 N7367 N7368 10
D7368 N7368 0 diode
R7369 N7368 N7369 10
D7369 N7369 0 diode
R7370 N7369 N7370 10
D7370 N7370 0 diode
R7371 N7370 N7371 10
D7371 N7371 0 diode
R7372 N7371 N7372 10
D7372 N7372 0 diode
R7373 N7372 N7373 10
D7373 N7373 0 diode
R7374 N7373 N7374 10
D7374 N7374 0 diode
R7375 N7374 N7375 10
D7375 N7375 0 diode
R7376 N7375 N7376 10
D7376 N7376 0 diode
R7377 N7376 N7377 10
D7377 N7377 0 diode
R7378 N7377 N7378 10
D7378 N7378 0 diode
R7379 N7378 N7379 10
D7379 N7379 0 diode
R7380 N7379 N7380 10
D7380 N7380 0 diode
R7381 N7380 N7381 10
D7381 N7381 0 diode
R7382 N7381 N7382 10
D7382 N7382 0 diode
R7383 N7382 N7383 10
D7383 N7383 0 diode
R7384 N7383 N7384 10
D7384 N7384 0 diode
R7385 N7384 N7385 10
D7385 N7385 0 diode
R7386 N7385 N7386 10
D7386 N7386 0 diode
R7387 N7386 N7387 10
D7387 N7387 0 diode
R7388 N7387 N7388 10
D7388 N7388 0 diode
R7389 N7388 N7389 10
D7389 N7389 0 diode
R7390 N7389 N7390 10
D7390 N7390 0 diode
R7391 N7390 N7391 10
D7391 N7391 0 diode
R7392 N7391 N7392 10
D7392 N7392 0 diode
R7393 N7392 N7393 10
D7393 N7393 0 diode
R7394 N7393 N7394 10
D7394 N7394 0 diode
R7395 N7394 N7395 10
D7395 N7395 0 diode
R7396 N7395 N7396 10
D7396 N7396 0 diode
R7397 N7396 N7397 10
D7397 N7397 0 diode
R7398 N7397 N7398 10
D7398 N7398 0 diode
R7399 N7398 N7399 10
D7399 N7399 0 diode
R7400 N7399 N7400 10
D7400 N7400 0 diode
R7401 N7400 N7401 10
D7401 N7401 0 diode
R7402 N7401 N7402 10
D7402 N7402 0 diode
R7403 N7402 N7403 10
D7403 N7403 0 diode
R7404 N7403 N7404 10
D7404 N7404 0 diode
R7405 N7404 N7405 10
D7405 N7405 0 diode
R7406 N7405 N7406 10
D7406 N7406 0 diode
R7407 N7406 N7407 10
D7407 N7407 0 diode
R7408 N7407 N7408 10
D7408 N7408 0 diode
R7409 N7408 N7409 10
D7409 N7409 0 diode
R7410 N7409 N7410 10
D7410 N7410 0 diode
R7411 N7410 N7411 10
D7411 N7411 0 diode
R7412 N7411 N7412 10
D7412 N7412 0 diode
R7413 N7412 N7413 10
D7413 N7413 0 diode
R7414 N7413 N7414 10
D7414 N7414 0 diode
R7415 N7414 N7415 10
D7415 N7415 0 diode
R7416 N7415 N7416 10
D7416 N7416 0 diode
R7417 N7416 N7417 10
D7417 N7417 0 diode
R7418 N7417 N7418 10
D7418 N7418 0 diode
R7419 N7418 N7419 10
D7419 N7419 0 diode
R7420 N7419 N7420 10
D7420 N7420 0 diode
R7421 N7420 N7421 10
D7421 N7421 0 diode
R7422 N7421 N7422 10
D7422 N7422 0 diode
R7423 N7422 N7423 10
D7423 N7423 0 diode
R7424 N7423 N7424 10
D7424 N7424 0 diode
R7425 N7424 N7425 10
D7425 N7425 0 diode
R7426 N7425 N7426 10
D7426 N7426 0 diode
R7427 N7426 N7427 10
D7427 N7427 0 diode
R7428 N7427 N7428 10
D7428 N7428 0 diode
R7429 N7428 N7429 10
D7429 N7429 0 diode
R7430 N7429 N7430 10
D7430 N7430 0 diode
R7431 N7430 N7431 10
D7431 N7431 0 diode
R7432 N7431 N7432 10
D7432 N7432 0 diode
R7433 N7432 N7433 10
D7433 N7433 0 diode
R7434 N7433 N7434 10
D7434 N7434 0 diode
R7435 N7434 N7435 10
D7435 N7435 0 diode
R7436 N7435 N7436 10
D7436 N7436 0 diode
R7437 N7436 N7437 10
D7437 N7437 0 diode
R7438 N7437 N7438 10
D7438 N7438 0 diode
R7439 N7438 N7439 10
D7439 N7439 0 diode
R7440 N7439 N7440 10
D7440 N7440 0 diode
R7441 N7440 N7441 10
D7441 N7441 0 diode
R7442 N7441 N7442 10
D7442 N7442 0 diode
R7443 N7442 N7443 10
D7443 N7443 0 diode
R7444 N7443 N7444 10
D7444 N7444 0 diode
R7445 N7444 N7445 10
D7445 N7445 0 diode
R7446 N7445 N7446 10
D7446 N7446 0 diode
R7447 N7446 N7447 10
D7447 N7447 0 diode
R7448 N7447 N7448 10
D7448 N7448 0 diode
R7449 N7448 N7449 10
D7449 N7449 0 diode
R7450 N7449 N7450 10
D7450 N7450 0 diode
R7451 N7450 N7451 10
D7451 N7451 0 diode
R7452 N7451 N7452 10
D7452 N7452 0 diode
R7453 N7452 N7453 10
D7453 N7453 0 diode
R7454 N7453 N7454 10
D7454 N7454 0 diode
R7455 N7454 N7455 10
D7455 N7455 0 diode
R7456 N7455 N7456 10
D7456 N7456 0 diode
R7457 N7456 N7457 10
D7457 N7457 0 diode
R7458 N7457 N7458 10
D7458 N7458 0 diode
R7459 N7458 N7459 10
D7459 N7459 0 diode
R7460 N7459 N7460 10
D7460 N7460 0 diode
R7461 N7460 N7461 10
D7461 N7461 0 diode
R7462 N7461 N7462 10
D7462 N7462 0 diode
R7463 N7462 N7463 10
D7463 N7463 0 diode
R7464 N7463 N7464 10
D7464 N7464 0 diode
R7465 N7464 N7465 10
D7465 N7465 0 diode
R7466 N7465 N7466 10
D7466 N7466 0 diode
R7467 N7466 N7467 10
D7467 N7467 0 diode
R7468 N7467 N7468 10
D7468 N7468 0 diode
R7469 N7468 N7469 10
D7469 N7469 0 diode
R7470 N7469 N7470 10
D7470 N7470 0 diode
R7471 N7470 N7471 10
D7471 N7471 0 diode
R7472 N7471 N7472 10
D7472 N7472 0 diode
R7473 N7472 N7473 10
D7473 N7473 0 diode
R7474 N7473 N7474 10
D7474 N7474 0 diode
R7475 N7474 N7475 10
D7475 N7475 0 diode
R7476 N7475 N7476 10
D7476 N7476 0 diode
R7477 N7476 N7477 10
D7477 N7477 0 diode
R7478 N7477 N7478 10
D7478 N7478 0 diode
R7479 N7478 N7479 10
D7479 N7479 0 diode
R7480 N7479 N7480 10
D7480 N7480 0 diode
R7481 N7480 N7481 10
D7481 N7481 0 diode
R7482 N7481 N7482 10
D7482 N7482 0 diode
R7483 N7482 N7483 10
D7483 N7483 0 diode
R7484 N7483 N7484 10
D7484 N7484 0 diode
R7485 N7484 N7485 10
D7485 N7485 0 diode
R7486 N7485 N7486 10
D7486 N7486 0 diode
R7487 N7486 N7487 10
D7487 N7487 0 diode
R7488 N7487 N7488 10
D7488 N7488 0 diode
R7489 N7488 N7489 10
D7489 N7489 0 diode
R7490 N7489 N7490 10
D7490 N7490 0 diode
R7491 N7490 N7491 10
D7491 N7491 0 diode
R7492 N7491 N7492 10
D7492 N7492 0 diode
R7493 N7492 N7493 10
D7493 N7493 0 diode
R7494 N7493 N7494 10
D7494 N7494 0 diode
R7495 N7494 N7495 10
D7495 N7495 0 diode
R7496 N7495 N7496 10
D7496 N7496 0 diode
R7497 N7496 N7497 10
D7497 N7497 0 diode
R7498 N7497 N7498 10
D7498 N7498 0 diode
R7499 N7498 N7499 10
D7499 N7499 0 diode
R7500 N7499 N7500 10
D7500 N7500 0 diode
R7501 N7500 N7501 10
D7501 N7501 0 diode
R7502 N7501 N7502 10
D7502 N7502 0 diode
R7503 N7502 N7503 10
D7503 N7503 0 diode
R7504 N7503 N7504 10
D7504 N7504 0 diode
R7505 N7504 N7505 10
D7505 N7505 0 diode
R7506 N7505 N7506 10
D7506 N7506 0 diode
R7507 N7506 N7507 10
D7507 N7507 0 diode
R7508 N7507 N7508 10
D7508 N7508 0 diode
R7509 N7508 N7509 10
D7509 N7509 0 diode
R7510 N7509 N7510 10
D7510 N7510 0 diode
R7511 N7510 N7511 10
D7511 N7511 0 diode
R7512 N7511 N7512 10
D7512 N7512 0 diode
R7513 N7512 N7513 10
D7513 N7513 0 diode
R7514 N7513 N7514 10
D7514 N7514 0 diode
R7515 N7514 N7515 10
D7515 N7515 0 diode
R7516 N7515 N7516 10
D7516 N7516 0 diode
R7517 N7516 N7517 10
D7517 N7517 0 diode
R7518 N7517 N7518 10
D7518 N7518 0 diode
R7519 N7518 N7519 10
D7519 N7519 0 diode
R7520 N7519 N7520 10
D7520 N7520 0 diode
R7521 N7520 N7521 10
D7521 N7521 0 diode
R7522 N7521 N7522 10
D7522 N7522 0 diode
R7523 N7522 N7523 10
D7523 N7523 0 diode
R7524 N7523 N7524 10
D7524 N7524 0 diode
R7525 N7524 N7525 10
D7525 N7525 0 diode
R7526 N7525 N7526 10
D7526 N7526 0 diode
R7527 N7526 N7527 10
D7527 N7527 0 diode
R7528 N7527 N7528 10
D7528 N7528 0 diode
R7529 N7528 N7529 10
D7529 N7529 0 diode
R7530 N7529 N7530 10
D7530 N7530 0 diode
R7531 N7530 N7531 10
D7531 N7531 0 diode
R7532 N7531 N7532 10
D7532 N7532 0 diode
R7533 N7532 N7533 10
D7533 N7533 0 diode
R7534 N7533 N7534 10
D7534 N7534 0 diode
R7535 N7534 N7535 10
D7535 N7535 0 diode
R7536 N7535 N7536 10
D7536 N7536 0 diode
R7537 N7536 N7537 10
D7537 N7537 0 diode
R7538 N7537 N7538 10
D7538 N7538 0 diode
R7539 N7538 N7539 10
D7539 N7539 0 diode
R7540 N7539 N7540 10
D7540 N7540 0 diode
R7541 N7540 N7541 10
D7541 N7541 0 diode
R7542 N7541 N7542 10
D7542 N7542 0 diode
R7543 N7542 N7543 10
D7543 N7543 0 diode
R7544 N7543 N7544 10
D7544 N7544 0 diode
R7545 N7544 N7545 10
D7545 N7545 0 diode
R7546 N7545 N7546 10
D7546 N7546 0 diode
R7547 N7546 N7547 10
D7547 N7547 0 diode
R7548 N7547 N7548 10
D7548 N7548 0 diode
R7549 N7548 N7549 10
D7549 N7549 0 diode
R7550 N7549 N7550 10
D7550 N7550 0 diode
R7551 N7550 N7551 10
D7551 N7551 0 diode
R7552 N7551 N7552 10
D7552 N7552 0 diode
R7553 N7552 N7553 10
D7553 N7553 0 diode
R7554 N7553 N7554 10
D7554 N7554 0 diode
R7555 N7554 N7555 10
D7555 N7555 0 diode
R7556 N7555 N7556 10
D7556 N7556 0 diode
R7557 N7556 N7557 10
D7557 N7557 0 diode
R7558 N7557 N7558 10
D7558 N7558 0 diode
R7559 N7558 N7559 10
D7559 N7559 0 diode
R7560 N7559 N7560 10
D7560 N7560 0 diode
R7561 N7560 N7561 10
D7561 N7561 0 diode
R7562 N7561 N7562 10
D7562 N7562 0 diode
R7563 N7562 N7563 10
D7563 N7563 0 diode
R7564 N7563 N7564 10
D7564 N7564 0 diode
R7565 N7564 N7565 10
D7565 N7565 0 diode
R7566 N7565 N7566 10
D7566 N7566 0 diode
R7567 N7566 N7567 10
D7567 N7567 0 diode
R7568 N7567 N7568 10
D7568 N7568 0 diode
R7569 N7568 N7569 10
D7569 N7569 0 diode
R7570 N7569 N7570 10
D7570 N7570 0 diode
R7571 N7570 N7571 10
D7571 N7571 0 diode
R7572 N7571 N7572 10
D7572 N7572 0 diode
R7573 N7572 N7573 10
D7573 N7573 0 diode
R7574 N7573 N7574 10
D7574 N7574 0 diode
R7575 N7574 N7575 10
D7575 N7575 0 diode
R7576 N7575 N7576 10
D7576 N7576 0 diode
R7577 N7576 N7577 10
D7577 N7577 0 diode
R7578 N7577 N7578 10
D7578 N7578 0 diode
R7579 N7578 N7579 10
D7579 N7579 0 diode
R7580 N7579 N7580 10
D7580 N7580 0 diode
R7581 N7580 N7581 10
D7581 N7581 0 diode
R7582 N7581 N7582 10
D7582 N7582 0 diode
R7583 N7582 N7583 10
D7583 N7583 0 diode
R7584 N7583 N7584 10
D7584 N7584 0 diode
R7585 N7584 N7585 10
D7585 N7585 0 diode
R7586 N7585 N7586 10
D7586 N7586 0 diode
R7587 N7586 N7587 10
D7587 N7587 0 diode
R7588 N7587 N7588 10
D7588 N7588 0 diode
R7589 N7588 N7589 10
D7589 N7589 0 diode
R7590 N7589 N7590 10
D7590 N7590 0 diode
R7591 N7590 N7591 10
D7591 N7591 0 diode
R7592 N7591 N7592 10
D7592 N7592 0 diode
R7593 N7592 N7593 10
D7593 N7593 0 diode
R7594 N7593 N7594 10
D7594 N7594 0 diode
R7595 N7594 N7595 10
D7595 N7595 0 diode
R7596 N7595 N7596 10
D7596 N7596 0 diode
R7597 N7596 N7597 10
D7597 N7597 0 diode
R7598 N7597 N7598 10
D7598 N7598 0 diode
R7599 N7598 N7599 10
D7599 N7599 0 diode
R7600 N7599 N7600 10
D7600 N7600 0 diode
R7601 N7600 N7601 10
D7601 N7601 0 diode
R7602 N7601 N7602 10
D7602 N7602 0 diode
R7603 N7602 N7603 10
D7603 N7603 0 diode
R7604 N7603 N7604 10
D7604 N7604 0 diode
R7605 N7604 N7605 10
D7605 N7605 0 diode
R7606 N7605 N7606 10
D7606 N7606 0 diode
R7607 N7606 N7607 10
D7607 N7607 0 diode
R7608 N7607 N7608 10
D7608 N7608 0 diode
R7609 N7608 N7609 10
D7609 N7609 0 diode
R7610 N7609 N7610 10
D7610 N7610 0 diode
R7611 N7610 N7611 10
D7611 N7611 0 diode
R7612 N7611 N7612 10
D7612 N7612 0 diode
R7613 N7612 N7613 10
D7613 N7613 0 diode
R7614 N7613 N7614 10
D7614 N7614 0 diode
R7615 N7614 N7615 10
D7615 N7615 0 diode
R7616 N7615 N7616 10
D7616 N7616 0 diode
R7617 N7616 N7617 10
D7617 N7617 0 diode
R7618 N7617 N7618 10
D7618 N7618 0 diode
R7619 N7618 N7619 10
D7619 N7619 0 diode
R7620 N7619 N7620 10
D7620 N7620 0 diode
R7621 N7620 N7621 10
D7621 N7621 0 diode
R7622 N7621 N7622 10
D7622 N7622 0 diode
R7623 N7622 N7623 10
D7623 N7623 0 diode
R7624 N7623 N7624 10
D7624 N7624 0 diode
R7625 N7624 N7625 10
D7625 N7625 0 diode
R7626 N7625 N7626 10
D7626 N7626 0 diode
R7627 N7626 N7627 10
D7627 N7627 0 diode
R7628 N7627 N7628 10
D7628 N7628 0 diode
R7629 N7628 N7629 10
D7629 N7629 0 diode
R7630 N7629 N7630 10
D7630 N7630 0 diode
R7631 N7630 N7631 10
D7631 N7631 0 diode
R7632 N7631 N7632 10
D7632 N7632 0 diode
R7633 N7632 N7633 10
D7633 N7633 0 diode
R7634 N7633 N7634 10
D7634 N7634 0 diode
R7635 N7634 N7635 10
D7635 N7635 0 diode
R7636 N7635 N7636 10
D7636 N7636 0 diode
R7637 N7636 N7637 10
D7637 N7637 0 diode
R7638 N7637 N7638 10
D7638 N7638 0 diode
R7639 N7638 N7639 10
D7639 N7639 0 diode
R7640 N7639 N7640 10
D7640 N7640 0 diode
R7641 N7640 N7641 10
D7641 N7641 0 diode
R7642 N7641 N7642 10
D7642 N7642 0 diode
R7643 N7642 N7643 10
D7643 N7643 0 diode
R7644 N7643 N7644 10
D7644 N7644 0 diode
R7645 N7644 N7645 10
D7645 N7645 0 diode
R7646 N7645 N7646 10
D7646 N7646 0 diode
R7647 N7646 N7647 10
D7647 N7647 0 diode
R7648 N7647 N7648 10
D7648 N7648 0 diode
R7649 N7648 N7649 10
D7649 N7649 0 diode
R7650 N7649 N7650 10
D7650 N7650 0 diode
R7651 N7650 N7651 10
D7651 N7651 0 diode
R7652 N7651 N7652 10
D7652 N7652 0 diode
R7653 N7652 N7653 10
D7653 N7653 0 diode
R7654 N7653 N7654 10
D7654 N7654 0 diode
R7655 N7654 N7655 10
D7655 N7655 0 diode
R7656 N7655 N7656 10
D7656 N7656 0 diode
R7657 N7656 N7657 10
D7657 N7657 0 diode
R7658 N7657 N7658 10
D7658 N7658 0 diode
R7659 N7658 N7659 10
D7659 N7659 0 diode
R7660 N7659 N7660 10
D7660 N7660 0 diode
R7661 N7660 N7661 10
D7661 N7661 0 diode
R7662 N7661 N7662 10
D7662 N7662 0 diode
R7663 N7662 N7663 10
D7663 N7663 0 diode
R7664 N7663 N7664 10
D7664 N7664 0 diode
R7665 N7664 N7665 10
D7665 N7665 0 diode
R7666 N7665 N7666 10
D7666 N7666 0 diode
R7667 N7666 N7667 10
D7667 N7667 0 diode
R7668 N7667 N7668 10
D7668 N7668 0 diode
R7669 N7668 N7669 10
D7669 N7669 0 diode
R7670 N7669 N7670 10
D7670 N7670 0 diode
R7671 N7670 N7671 10
D7671 N7671 0 diode
R7672 N7671 N7672 10
D7672 N7672 0 diode
R7673 N7672 N7673 10
D7673 N7673 0 diode
R7674 N7673 N7674 10
D7674 N7674 0 diode
R7675 N7674 N7675 10
D7675 N7675 0 diode
R7676 N7675 N7676 10
D7676 N7676 0 diode
R7677 N7676 N7677 10
D7677 N7677 0 diode
R7678 N7677 N7678 10
D7678 N7678 0 diode
R7679 N7678 N7679 10
D7679 N7679 0 diode
R7680 N7679 N7680 10
D7680 N7680 0 diode
R7681 N7680 N7681 10
D7681 N7681 0 diode
R7682 N7681 N7682 10
D7682 N7682 0 diode
R7683 N7682 N7683 10
D7683 N7683 0 diode
R7684 N7683 N7684 10
D7684 N7684 0 diode
R7685 N7684 N7685 10
D7685 N7685 0 diode
R7686 N7685 N7686 10
D7686 N7686 0 diode
R7687 N7686 N7687 10
D7687 N7687 0 diode
R7688 N7687 N7688 10
D7688 N7688 0 diode
R7689 N7688 N7689 10
D7689 N7689 0 diode
R7690 N7689 N7690 10
D7690 N7690 0 diode
R7691 N7690 N7691 10
D7691 N7691 0 diode
R7692 N7691 N7692 10
D7692 N7692 0 diode
R7693 N7692 N7693 10
D7693 N7693 0 diode
R7694 N7693 N7694 10
D7694 N7694 0 diode
R7695 N7694 N7695 10
D7695 N7695 0 diode
R7696 N7695 N7696 10
D7696 N7696 0 diode
R7697 N7696 N7697 10
D7697 N7697 0 diode
R7698 N7697 N7698 10
D7698 N7698 0 diode
R7699 N7698 N7699 10
D7699 N7699 0 diode
R7700 N7699 N7700 10
D7700 N7700 0 diode
R7701 N7700 N7701 10
D7701 N7701 0 diode
R7702 N7701 N7702 10
D7702 N7702 0 diode
R7703 N7702 N7703 10
D7703 N7703 0 diode
R7704 N7703 N7704 10
D7704 N7704 0 diode
R7705 N7704 N7705 10
D7705 N7705 0 diode
R7706 N7705 N7706 10
D7706 N7706 0 diode
R7707 N7706 N7707 10
D7707 N7707 0 diode
R7708 N7707 N7708 10
D7708 N7708 0 diode
R7709 N7708 N7709 10
D7709 N7709 0 diode
R7710 N7709 N7710 10
D7710 N7710 0 diode
R7711 N7710 N7711 10
D7711 N7711 0 diode
R7712 N7711 N7712 10
D7712 N7712 0 diode
R7713 N7712 N7713 10
D7713 N7713 0 diode
R7714 N7713 N7714 10
D7714 N7714 0 diode
R7715 N7714 N7715 10
D7715 N7715 0 diode
R7716 N7715 N7716 10
D7716 N7716 0 diode
R7717 N7716 N7717 10
D7717 N7717 0 diode
R7718 N7717 N7718 10
D7718 N7718 0 diode
R7719 N7718 N7719 10
D7719 N7719 0 diode
R7720 N7719 N7720 10
D7720 N7720 0 diode
R7721 N7720 N7721 10
D7721 N7721 0 diode
R7722 N7721 N7722 10
D7722 N7722 0 diode
R7723 N7722 N7723 10
D7723 N7723 0 diode
R7724 N7723 N7724 10
D7724 N7724 0 diode
R7725 N7724 N7725 10
D7725 N7725 0 diode
R7726 N7725 N7726 10
D7726 N7726 0 diode
R7727 N7726 N7727 10
D7727 N7727 0 diode
R7728 N7727 N7728 10
D7728 N7728 0 diode
R7729 N7728 N7729 10
D7729 N7729 0 diode
R7730 N7729 N7730 10
D7730 N7730 0 diode
R7731 N7730 N7731 10
D7731 N7731 0 diode
R7732 N7731 N7732 10
D7732 N7732 0 diode
R7733 N7732 N7733 10
D7733 N7733 0 diode
R7734 N7733 N7734 10
D7734 N7734 0 diode
R7735 N7734 N7735 10
D7735 N7735 0 diode
R7736 N7735 N7736 10
D7736 N7736 0 diode
R7737 N7736 N7737 10
D7737 N7737 0 diode
R7738 N7737 N7738 10
D7738 N7738 0 diode
R7739 N7738 N7739 10
D7739 N7739 0 diode
R7740 N7739 N7740 10
D7740 N7740 0 diode
R7741 N7740 N7741 10
D7741 N7741 0 diode
R7742 N7741 N7742 10
D7742 N7742 0 diode
R7743 N7742 N7743 10
D7743 N7743 0 diode
R7744 N7743 N7744 10
D7744 N7744 0 diode
R7745 N7744 N7745 10
D7745 N7745 0 diode
R7746 N7745 N7746 10
D7746 N7746 0 diode
R7747 N7746 N7747 10
D7747 N7747 0 diode
R7748 N7747 N7748 10
D7748 N7748 0 diode
R7749 N7748 N7749 10
D7749 N7749 0 diode
R7750 N7749 N7750 10
D7750 N7750 0 diode
R7751 N7750 N7751 10
D7751 N7751 0 diode
R7752 N7751 N7752 10
D7752 N7752 0 diode
R7753 N7752 N7753 10
D7753 N7753 0 diode
R7754 N7753 N7754 10
D7754 N7754 0 diode
R7755 N7754 N7755 10
D7755 N7755 0 diode
R7756 N7755 N7756 10
D7756 N7756 0 diode
R7757 N7756 N7757 10
D7757 N7757 0 diode
R7758 N7757 N7758 10
D7758 N7758 0 diode
R7759 N7758 N7759 10
D7759 N7759 0 diode
R7760 N7759 N7760 10
D7760 N7760 0 diode
R7761 N7760 N7761 10
D7761 N7761 0 diode
R7762 N7761 N7762 10
D7762 N7762 0 diode
R7763 N7762 N7763 10
D7763 N7763 0 diode
R7764 N7763 N7764 10
D7764 N7764 0 diode
R7765 N7764 N7765 10
D7765 N7765 0 diode
R7766 N7765 N7766 10
D7766 N7766 0 diode
R7767 N7766 N7767 10
D7767 N7767 0 diode
R7768 N7767 N7768 10
D7768 N7768 0 diode
R7769 N7768 N7769 10
D7769 N7769 0 diode
R7770 N7769 N7770 10
D7770 N7770 0 diode
R7771 N7770 N7771 10
D7771 N7771 0 diode
R7772 N7771 N7772 10
D7772 N7772 0 diode
R7773 N7772 N7773 10
D7773 N7773 0 diode
R7774 N7773 N7774 10
D7774 N7774 0 diode
R7775 N7774 N7775 10
D7775 N7775 0 diode
R7776 N7775 N7776 10
D7776 N7776 0 diode
R7777 N7776 N7777 10
D7777 N7777 0 diode
R7778 N7777 N7778 10
D7778 N7778 0 diode
R7779 N7778 N7779 10
D7779 N7779 0 diode
R7780 N7779 N7780 10
D7780 N7780 0 diode
R7781 N7780 N7781 10
D7781 N7781 0 diode
R7782 N7781 N7782 10
D7782 N7782 0 diode
R7783 N7782 N7783 10
D7783 N7783 0 diode
R7784 N7783 N7784 10
D7784 N7784 0 diode
R7785 N7784 N7785 10
D7785 N7785 0 diode
R7786 N7785 N7786 10
D7786 N7786 0 diode
R7787 N7786 N7787 10
D7787 N7787 0 diode
R7788 N7787 N7788 10
D7788 N7788 0 diode
R7789 N7788 N7789 10
D7789 N7789 0 diode
R7790 N7789 N7790 10
D7790 N7790 0 diode
R7791 N7790 N7791 10
D7791 N7791 0 diode
R7792 N7791 N7792 10
D7792 N7792 0 diode
R7793 N7792 N7793 10
D7793 N7793 0 diode
R7794 N7793 N7794 10
D7794 N7794 0 diode
R7795 N7794 N7795 10
D7795 N7795 0 diode
R7796 N7795 N7796 10
D7796 N7796 0 diode
R7797 N7796 N7797 10
D7797 N7797 0 diode
R7798 N7797 N7798 10
D7798 N7798 0 diode
R7799 N7798 N7799 10
D7799 N7799 0 diode
R7800 N7799 N7800 10
D7800 N7800 0 diode
R7801 N7800 N7801 10
D7801 N7801 0 diode
R7802 N7801 N7802 10
D7802 N7802 0 diode
R7803 N7802 N7803 10
D7803 N7803 0 diode
R7804 N7803 N7804 10
D7804 N7804 0 diode
R7805 N7804 N7805 10
D7805 N7805 0 diode
R7806 N7805 N7806 10
D7806 N7806 0 diode
R7807 N7806 N7807 10
D7807 N7807 0 diode
R7808 N7807 N7808 10
D7808 N7808 0 diode
R7809 N7808 N7809 10
D7809 N7809 0 diode
R7810 N7809 N7810 10
D7810 N7810 0 diode
R7811 N7810 N7811 10
D7811 N7811 0 diode
R7812 N7811 N7812 10
D7812 N7812 0 diode
R7813 N7812 N7813 10
D7813 N7813 0 diode
R7814 N7813 N7814 10
D7814 N7814 0 diode
R7815 N7814 N7815 10
D7815 N7815 0 diode
R7816 N7815 N7816 10
D7816 N7816 0 diode
R7817 N7816 N7817 10
D7817 N7817 0 diode
R7818 N7817 N7818 10
D7818 N7818 0 diode
R7819 N7818 N7819 10
D7819 N7819 0 diode
R7820 N7819 N7820 10
D7820 N7820 0 diode
R7821 N7820 N7821 10
D7821 N7821 0 diode
R7822 N7821 N7822 10
D7822 N7822 0 diode
R7823 N7822 N7823 10
D7823 N7823 0 diode
R7824 N7823 N7824 10
D7824 N7824 0 diode
R7825 N7824 N7825 10
D7825 N7825 0 diode
R7826 N7825 N7826 10
D7826 N7826 0 diode
R7827 N7826 N7827 10
D7827 N7827 0 diode
R7828 N7827 N7828 10
D7828 N7828 0 diode
R7829 N7828 N7829 10
D7829 N7829 0 diode
R7830 N7829 N7830 10
D7830 N7830 0 diode
R7831 N7830 N7831 10
D7831 N7831 0 diode
R7832 N7831 N7832 10
D7832 N7832 0 diode
R7833 N7832 N7833 10
D7833 N7833 0 diode
R7834 N7833 N7834 10
D7834 N7834 0 diode
R7835 N7834 N7835 10
D7835 N7835 0 diode
R7836 N7835 N7836 10
D7836 N7836 0 diode
R7837 N7836 N7837 10
D7837 N7837 0 diode
R7838 N7837 N7838 10
D7838 N7838 0 diode
R7839 N7838 N7839 10
D7839 N7839 0 diode
R7840 N7839 N7840 10
D7840 N7840 0 diode
R7841 N7840 N7841 10
D7841 N7841 0 diode
R7842 N7841 N7842 10
D7842 N7842 0 diode
R7843 N7842 N7843 10
D7843 N7843 0 diode
R7844 N7843 N7844 10
D7844 N7844 0 diode
R7845 N7844 N7845 10
D7845 N7845 0 diode
R7846 N7845 N7846 10
D7846 N7846 0 diode
R7847 N7846 N7847 10
D7847 N7847 0 diode
R7848 N7847 N7848 10
D7848 N7848 0 diode
R7849 N7848 N7849 10
D7849 N7849 0 diode
R7850 N7849 N7850 10
D7850 N7850 0 diode
R7851 N7850 N7851 10
D7851 N7851 0 diode
R7852 N7851 N7852 10
D7852 N7852 0 diode
R7853 N7852 N7853 10
D7853 N7853 0 diode
R7854 N7853 N7854 10
D7854 N7854 0 diode
R7855 N7854 N7855 10
D7855 N7855 0 diode
R7856 N7855 N7856 10
D7856 N7856 0 diode
R7857 N7856 N7857 10
D7857 N7857 0 diode
R7858 N7857 N7858 10
D7858 N7858 0 diode
R7859 N7858 N7859 10
D7859 N7859 0 diode
R7860 N7859 N7860 10
D7860 N7860 0 diode
R7861 N7860 N7861 10
D7861 N7861 0 diode
R7862 N7861 N7862 10
D7862 N7862 0 diode
R7863 N7862 N7863 10
D7863 N7863 0 diode
R7864 N7863 N7864 10
D7864 N7864 0 diode
R7865 N7864 N7865 10
D7865 N7865 0 diode
R7866 N7865 N7866 10
D7866 N7866 0 diode
R7867 N7866 N7867 10
D7867 N7867 0 diode
R7868 N7867 N7868 10
D7868 N7868 0 diode
R7869 N7868 N7869 10
D7869 N7869 0 diode
R7870 N7869 N7870 10
D7870 N7870 0 diode
R7871 N7870 N7871 10
D7871 N7871 0 diode
R7872 N7871 N7872 10
D7872 N7872 0 diode
R7873 N7872 N7873 10
D7873 N7873 0 diode
R7874 N7873 N7874 10
D7874 N7874 0 diode
R7875 N7874 N7875 10
D7875 N7875 0 diode
R7876 N7875 N7876 10
D7876 N7876 0 diode
R7877 N7876 N7877 10
D7877 N7877 0 diode
R7878 N7877 N7878 10
D7878 N7878 0 diode
R7879 N7878 N7879 10
D7879 N7879 0 diode
R7880 N7879 N7880 10
D7880 N7880 0 diode
R7881 N7880 N7881 10
D7881 N7881 0 diode
R7882 N7881 N7882 10
D7882 N7882 0 diode
R7883 N7882 N7883 10
D7883 N7883 0 diode
R7884 N7883 N7884 10
D7884 N7884 0 diode
R7885 N7884 N7885 10
D7885 N7885 0 diode
R7886 N7885 N7886 10
D7886 N7886 0 diode
R7887 N7886 N7887 10
D7887 N7887 0 diode
R7888 N7887 N7888 10
D7888 N7888 0 diode
R7889 N7888 N7889 10
D7889 N7889 0 diode
R7890 N7889 N7890 10
D7890 N7890 0 diode
R7891 N7890 N7891 10
D7891 N7891 0 diode
R7892 N7891 N7892 10
D7892 N7892 0 diode
R7893 N7892 N7893 10
D7893 N7893 0 diode
R7894 N7893 N7894 10
D7894 N7894 0 diode
R7895 N7894 N7895 10
D7895 N7895 0 diode
R7896 N7895 N7896 10
D7896 N7896 0 diode
R7897 N7896 N7897 10
D7897 N7897 0 diode
R7898 N7897 N7898 10
D7898 N7898 0 diode
R7899 N7898 N7899 10
D7899 N7899 0 diode
R7900 N7899 N7900 10
D7900 N7900 0 diode
R7901 N7900 N7901 10
D7901 N7901 0 diode
R7902 N7901 N7902 10
D7902 N7902 0 diode
R7903 N7902 N7903 10
D7903 N7903 0 diode
R7904 N7903 N7904 10
D7904 N7904 0 diode
R7905 N7904 N7905 10
D7905 N7905 0 diode
R7906 N7905 N7906 10
D7906 N7906 0 diode
R7907 N7906 N7907 10
D7907 N7907 0 diode
R7908 N7907 N7908 10
D7908 N7908 0 diode
R7909 N7908 N7909 10
D7909 N7909 0 diode
R7910 N7909 N7910 10
D7910 N7910 0 diode
R7911 N7910 N7911 10
D7911 N7911 0 diode
R7912 N7911 N7912 10
D7912 N7912 0 diode
R7913 N7912 N7913 10
D7913 N7913 0 diode
R7914 N7913 N7914 10
D7914 N7914 0 diode
R7915 N7914 N7915 10
D7915 N7915 0 diode
R7916 N7915 N7916 10
D7916 N7916 0 diode
R7917 N7916 N7917 10
D7917 N7917 0 diode
R7918 N7917 N7918 10
D7918 N7918 0 diode
R7919 N7918 N7919 10
D7919 N7919 0 diode
R7920 N7919 N7920 10
D7920 N7920 0 diode
R7921 N7920 N7921 10
D7921 N7921 0 diode
R7922 N7921 N7922 10
D7922 N7922 0 diode
R7923 N7922 N7923 10
D7923 N7923 0 diode
R7924 N7923 N7924 10
D7924 N7924 0 diode
R7925 N7924 N7925 10
D7925 N7925 0 diode
R7926 N7925 N7926 10
D7926 N7926 0 diode
R7927 N7926 N7927 10
D7927 N7927 0 diode
R7928 N7927 N7928 10
D7928 N7928 0 diode
R7929 N7928 N7929 10
D7929 N7929 0 diode
R7930 N7929 N7930 10
D7930 N7930 0 diode
R7931 N7930 N7931 10
D7931 N7931 0 diode
R7932 N7931 N7932 10
D7932 N7932 0 diode
R7933 N7932 N7933 10
D7933 N7933 0 diode
R7934 N7933 N7934 10
D7934 N7934 0 diode
R7935 N7934 N7935 10
D7935 N7935 0 diode
R7936 N7935 N7936 10
D7936 N7936 0 diode
R7937 N7936 N7937 10
D7937 N7937 0 diode
R7938 N7937 N7938 10
D7938 N7938 0 diode
R7939 N7938 N7939 10
D7939 N7939 0 diode
R7940 N7939 N7940 10
D7940 N7940 0 diode
R7941 N7940 N7941 10
D7941 N7941 0 diode
R7942 N7941 N7942 10
D7942 N7942 0 diode
R7943 N7942 N7943 10
D7943 N7943 0 diode
R7944 N7943 N7944 10
D7944 N7944 0 diode
R7945 N7944 N7945 10
D7945 N7945 0 diode
R7946 N7945 N7946 10
D7946 N7946 0 diode
R7947 N7946 N7947 10
D7947 N7947 0 diode
R7948 N7947 N7948 10
D7948 N7948 0 diode
R7949 N7948 N7949 10
D7949 N7949 0 diode
R7950 N7949 N7950 10
D7950 N7950 0 diode
R7951 N7950 N7951 10
D7951 N7951 0 diode
R7952 N7951 N7952 10
D7952 N7952 0 diode
R7953 N7952 N7953 10
D7953 N7953 0 diode
R7954 N7953 N7954 10
D7954 N7954 0 diode
R7955 N7954 N7955 10
D7955 N7955 0 diode
R7956 N7955 N7956 10
D7956 N7956 0 diode
R7957 N7956 N7957 10
D7957 N7957 0 diode
R7958 N7957 N7958 10
D7958 N7958 0 diode
R7959 N7958 N7959 10
D7959 N7959 0 diode
R7960 N7959 N7960 10
D7960 N7960 0 diode
R7961 N7960 N7961 10
D7961 N7961 0 diode
R7962 N7961 N7962 10
D7962 N7962 0 diode
R7963 N7962 N7963 10
D7963 N7963 0 diode
R7964 N7963 N7964 10
D7964 N7964 0 diode
R7965 N7964 N7965 10
D7965 N7965 0 diode
R7966 N7965 N7966 10
D7966 N7966 0 diode
R7967 N7966 N7967 10
D7967 N7967 0 diode
R7968 N7967 N7968 10
D7968 N7968 0 diode
R7969 N7968 N7969 10
D7969 N7969 0 diode
R7970 N7969 N7970 10
D7970 N7970 0 diode
R7971 N7970 N7971 10
D7971 N7971 0 diode
R7972 N7971 N7972 10
D7972 N7972 0 diode
R7973 N7972 N7973 10
D7973 N7973 0 diode
R7974 N7973 N7974 10
D7974 N7974 0 diode
R7975 N7974 N7975 10
D7975 N7975 0 diode
R7976 N7975 N7976 10
D7976 N7976 0 diode
R7977 N7976 N7977 10
D7977 N7977 0 diode
R7978 N7977 N7978 10
D7978 N7978 0 diode
R7979 N7978 N7979 10
D7979 N7979 0 diode
R7980 N7979 N7980 10
D7980 N7980 0 diode
R7981 N7980 N7981 10
D7981 N7981 0 diode
R7982 N7981 N7982 10
D7982 N7982 0 diode
R7983 N7982 N7983 10
D7983 N7983 0 diode
R7984 N7983 N7984 10
D7984 N7984 0 diode
R7985 N7984 N7985 10
D7985 N7985 0 diode
R7986 N7985 N7986 10
D7986 N7986 0 diode
R7987 N7986 N7987 10
D7987 N7987 0 diode
R7988 N7987 N7988 10
D7988 N7988 0 diode
R7989 N7988 N7989 10
D7989 N7989 0 diode
R7990 N7989 N7990 10
D7990 N7990 0 diode
R7991 N7990 N7991 10
D7991 N7991 0 diode
R7992 N7991 N7992 10
D7992 N7992 0 diode
R7993 N7992 N7993 10
D7993 N7993 0 diode
R7994 N7993 N7994 10
D7994 N7994 0 diode
R7995 N7994 N7995 10
D7995 N7995 0 diode
R7996 N7995 N7996 10
D7996 N7996 0 diode
R7997 N7996 N7997 10
D7997 N7997 0 diode
R7998 N7997 N7998 10
D7998 N7998 0 diode
R7999 N7998 N7999 10
D7999 N7999 0 diode
R8000 N7999 N8000 10
D8000 N8000 0 diode
R8001 N8000 N8001 10
D8001 N8001 0 diode
R8002 N8001 N8002 10
D8002 N8002 0 diode
R8003 N8002 N8003 10
D8003 N8003 0 diode
R8004 N8003 N8004 10
D8004 N8004 0 diode
R8005 N8004 N8005 10
D8005 N8005 0 diode
R8006 N8005 N8006 10
D8006 N8006 0 diode
R8007 N8006 N8007 10
D8007 N8007 0 diode
R8008 N8007 N8008 10
D8008 N8008 0 diode
R8009 N8008 N8009 10
D8009 N8009 0 diode
R8010 N8009 N8010 10
D8010 N8010 0 diode
R8011 N8010 N8011 10
D8011 N8011 0 diode
R8012 N8011 N8012 10
D8012 N8012 0 diode
R8013 N8012 N8013 10
D8013 N8013 0 diode
R8014 N8013 N8014 10
D8014 N8014 0 diode
R8015 N8014 N8015 10
D8015 N8015 0 diode
R8016 N8015 N8016 10
D8016 N8016 0 diode
R8017 N8016 N8017 10
D8017 N8017 0 diode
R8018 N8017 N8018 10
D8018 N8018 0 diode
R8019 N8018 N8019 10
D8019 N8019 0 diode
R8020 N8019 N8020 10
D8020 N8020 0 diode
R8021 N8020 N8021 10
D8021 N8021 0 diode
R8022 N8021 N8022 10
D8022 N8022 0 diode
R8023 N8022 N8023 10
D8023 N8023 0 diode
R8024 N8023 N8024 10
D8024 N8024 0 diode
R8025 N8024 N8025 10
D8025 N8025 0 diode
R8026 N8025 N8026 10
D8026 N8026 0 diode
R8027 N8026 N8027 10
D8027 N8027 0 diode
R8028 N8027 N8028 10
D8028 N8028 0 diode
R8029 N8028 N8029 10
D8029 N8029 0 diode
R8030 N8029 N8030 10
D8030 N8030 0 diode
R8031 N8030 N8031 10
D8031 N8031 0 diode
R8032 N8031 N8032 10
D8032 N8032 0 diode
R8033 N8032 N8033 10
D8033 N8033 0 diode
R8034 N8033 N8034 10
D8034 N8034 0 diode
R8035 N8034 N8035 10
D8035 N8035 0 diode
R8036 N8035 N8036 10
D8036 N8036 0 diode
R8037 N8036 N8037 10
D8037 N8037 0 diode
R8038 N8037 N8038 10
D8038 N8038 0 diode
R8039 N8038 N8039 10
D8039 N8039 0 diode
R8040 N8039 N8040 10
D8040 N8040 0 diode
R8041 N8040 N8041 10
D8041 N8041 0 diode
R8042 N8041 N8042 10
D8042 N8042 0 diode
R8043 N8042 N8043 10
D8043 N8043 0 diode
R8044 N8043 N8044 10
D8044 N8044 0 diode
R8045 N8044 N8045 10
D8045 N8045 0 diode
R8046 N8045 N8046 10
D8046 N8046 0 diode
R8047 N8046 N8047 10
D8047 N8047 0 diode
R8048 N8047 N8048 10
D8048 N8048 0 diode
R8049 N8048 N8049 10
D8049 N8049 0 diode
R8050 N8049 N8050 10
D8050 N8050 0 diode
R8051 N8050 N8051 10
D8051 N8051 0 diode
R8052 N8051 N8052 10
D8052 N8052 0 diode
R8053 N8052 N8053 10
D8053 N8053 0 diode
R8054 N8053 N8054 10
D8054 N8054 0 diode
R8055 N8054 N8055 10
D8055 N8055 0 diode
R8056 N8055 N8056 10
D8056 N8056 0 diode
R8057 N8056 N8057 10
D8057 N8057 0 diode
R8058 N8057 N8058 10
D8058 N8058 0 diode
R8059 N8058 N8059 10
D8059 N8059 0 diode
R8060 N8059 N8060 10
D8060 N8060 0 diode
R8061 N8060 N8061 10
D8061 N8061 0 diode
R8062 N8061 N8062 10
D8062 N8062 0 diode
R8063 N8062 N8063 10
D8063 N8063 0 diode
R8064 N8063 N8064 10
D8064 N8064 0 diode
R8065 N8064 N8065 10
D8065 N8065 0 diode
R8066 N8065 N8066 10
D8066 N8066 0 diode
R8067 N8066 N8067 10
D8067 N8067 0 diode
R8068 N8067 N8068 10
D8068 N8068 0 diode
R8069 N8068 N8069 10
D8069 N8069 0 diode
R8070 N8069 N8070 10
D8070 N8070 0 diode
R8071 N8070 N8071 10
D8071 N8071 0 diode
R8072 N8071 N8072 10
D8072 N8072 0 diode
R8073 N8072 N8073 10
D8073 N8073 0 diode
R8074 N8073 N8074 10
D8074 N8074 0 diode
R8075 N8074 N8075 10
D8075 N8075 0 diode
R8076 N8075 N8076 10
D8076 N8076 0 diode
R8077 N8076 N8077 10
D8077 N8077 0 diode
R8078 N8077 N8078 10
D8078 N8078 0 diode
R8079 N8078 N8079 10
D8079 N8079 0 diode
R8080 N8079 N8080 10
D8080 N8080 0 diode
R8081 N8080 N8081 10
D8081 N8081 0 diode
R8082 N8081 N8082 10
D8082 N8082 0 diode
R8083 N8082 N8083 10
D8083 N8083 0 diode
R8084 N8083 N8084 10
D8084 N8084 0 diode
R8085 N8084 N8085 10
D8085 N8085 0 diode
R8086 N8085 N8086 10
D8086 N8086 0 diode
R8087 N8086 N8087 10
D8087 N8087 0 diode
R8088 N8087 N8088 10
D8088 N8088 0 diode
R8089 N8088 N8089 10
D8089 N8089 0 diode
R8090 N8089 N8090 10
D8090 N8090 0 diode
R8091 N8090 N8091 10
D8091 N8091 0 diode
R8092 N8091 N8092 10
D8092 N8092 0 diode
R8093 N8092 N8093 10
D8093 N8093 0 diode
R8094 N8093 N8094 10
D8094 N8094 0 diode
R8095 N8094 N8095 10
D8095 N8095 0 diode
R8096 N8095 N8096 10
D8096 N8096 0 diode
R8097 N8096 N8097 10
D8097 N8097 0 diode
R8098 N8097 N8098 10
D8098 N8098 0 diode
R8099 N8098 N8099 10
D8099 N8099 0 diode
R8100 N8099 N8100 10
D8100 N8100 0 diode
R8101 N8100 N8101 10
D8101 N8101 0 diode
R8102 N8101 N8102 10
D8102 N8102 0 diode
R8103 N8102 N8103 10
D8103 N8103 0 diode
R8104 N8103 N8104 10
D8104 N8104 0 diode
R8105 N8104 N8105 10
D8105 N8105 0 diode
R8106 N8105 N8106 10
D8106 N8106 0 diode
R8107 N8106 N8107 10
D8107 N8107 0 diode
R8108 N8107 N8108 10
D8108 N8108 0 diode
R8109 N8108 N8109 10
D8109 N8109 0 diode
R8110 N8109 N8110 10
D8110 N8110 0 diode
R8111 N8110 N8111 10
D8111 N8111 0 diode
R8112 N8111 N8112 10
D8112 N8112 0 diode
R8113 N8112 N8113 10
D8113 N8113 0 diode
R8114 N8113 N8114 10
D8114 N8114 0 diode
R8115 N8114 N8115 10
D8115 N8115 0 diode
R8116 N8115 N8116 10
D8116 N8116 0 diode
R8117 N8116 N8117 10
D8117 N8117 0 diode
R8118 N8117 N8118 10
D8118 N8118 0 diode
R8119 N8118 N8119 10
D8119 N8119 0 diode
R8120 N8119 N8120 10
D8120 N8120 0 diode
R8121 N8120 N8121 10
D8121 N8121 0 diode
R8122 N8121 N8122 10
D8122 N8122 0 diode
R8123 N8122 N8123 10
D8123 N8123 0 diode
R8124 N8123 N8124 10
D8124 N8124 0 diode
R8125 N8124 N8125 10
D8125 N8125 0 diode
R8126 N8125 N8126 10
D8126 N8126 0 diode
R8127 N8126 N8127 10
D8127 N8127 0 diode
R8128 N8127 N8128 10
D8128 N8128 0 diode
R8129 N8128 N8129 10
D8129 N8129 0 diode
R8130 N8129 N8130 10
D8130 N8130 0 diode
R8131 N8130 N8131 10
D8131 N8131 0 diode
R8132 N8131 N8132 10
D8132 N8132 0 diode
R8133 N8132 N8133 10
D8133 N8133 0 diode
R8134 N8133 N8134 10
D8134 N8134 0 diode
R8135 N8134 N8135 10
D8135 N8135 0 diode
R8136 N8135 N8136 10
D8136 N8136 0 diode
R8137 N8136 N8137 10
D8137 N8137 0 diode
R8138 N8137 N8138 10
D8138 N8138 0 diode
R8139 N8138 N8139 10
D8139 N8139 0 diode
R8140 N8139 N8140 10
D8140 N8140 0 diode
R8141 N8140 N8141 10
D8141 N8141 0 diode
R8142 N8141 N8142 10
D8142 N8142 0 diode
R8143 N8142 N8143 10
D8143 N8143 0 diode
R8144 N8143 N8144 10
D8144 N8144 0 diode
R8145 N8144 N8145 10
D8145 N8145 0 diode
R8146 N8145 N8146 10
D8146 N8146 0 diode
R8147 N8146 N8147 10
D8147 N8147 0 diode
R8148 N8147 N8148 10
D8148 N8148 0 diode
R8149 N8148 N8149 10
D8149 N8149 0 diode
R8150 N8149 N8150 10
D8150 N8150 0 diode
R8151 N8150 N8151 10
D8151 N8151 0 diode
R8152 N8151 N8152 10
D8152 N8152 0 diode
R8153 N8152 N8153 10
D8153 N8153 0 diode
R8154 N8153 N8154 10
D8154 N8154 0 diode
R8155 N8154 N8155 10
D8155 N8155 0 diode
R8156 N8155 N8156 10
D8156 N8156 0 diode
R8157 N8156 N8157 10
D8157 N8157 0 diode
R8158 N8157 N8158 10
D8158 N8158 0 diode
R8159 N8158 N8159 10
D8159 N8159 0 diode
R8160 N8159 N8160 10
D8160 N8160 0 diode
R8161 N8160 N8161 10
D8161 N8161 0 diode
R8162 N8161 N8162 10
D8162 N8162 0 diode
R8163 N8162 N8163 10
D8163 N8163 0 diode
R8164 N8163 N8164 10
D8164 N8164 0 diode
R8165 N8164 N8165 10
D8165 N8165 0 diode
R8166 N8165 N8166 10
D8166 N8166 0 diode
R8167 N8166 N8167 10
D8167 N8167 0 diode
R8168 N8167 N8168 10
D8168 N8168 0 diode
R8169 N8168 N8169 10
D8169 N8169 0 diode
R8170 N8169 N8170 10
D8170 N8170 0 diode
R8171 N8170 N8171 10
D8171 N8171 0 diode
R8172 N8171 N8172 10
D8172 N8172 0 diode
R8173 N8172 N8173 10
D8173 N8173 0 diode
R8174 N8173 N8174 10
D8174 N8174 0 diode
R8175 N8174 N8175 10
D8175 N8175 0 diode
R8176 N8175 N8176 10
D8176 N8176 0 diode
R8177 N8176 N8177 10
D8177 N8177 0 diode
R8178 N8177 N8178 10
D8178 N8178 0 diode
R8179 N8178 N8179 10
D8179 N8179 0 diode
R8180 N8179 N8180 10
D8180 N8180 0 diode
R8181 N8180 N8181 10
D8181 N8181 0 diode
R8182 N8181 N8182 10
D8182 N8182 0 diode
R8183 N8182 N8183 10
D8183 N8183 0 diode
R8184 N8183 N8184 10
D8184 N8184 0 diode
R8185 N8184 N8185 10
D8185 N8185 0 diode
R8186 N8185 N8186 10
D8186 N8186 0 diode
R8187 N8186 N8187 10
D8187 N8187 0 diode
R8188 N8187 N8188 10
D8188 N8188 0 diode
R8189 N8188 N8189 10
D8189 N8189 0 diode
R8190 N8189 N8190 10
D8190 N8190 0 diode
R8191 N8190 N8191 10
D8191 N8191 0 diode
R8192 N8191 N8192 10
D8192 N8192 0 diode
R8193 N8192 N8193 10
D8193 N8193 0 diode
R8194 N8193 N8194 10
D8194 N8194 0 diode
R8195 N8194 N8195 10
D8195 N8195 0 diode
R8196 N8195 N8196 10
D8196 N8196 0 diode
R8197 N8196 N8197 10
D8197 N8197 0 diode
R8198 N8197 N8198 10
D8198 N8198 0 diode
R8199 N8198 N8199 10
D8199 N8199 0 diode
R8200 N8199 N8200 10
D8200 N8200 0 diode
R8201 N8200 N8201 10
D8201 N8201 0 diode
R8202 N8201 N8202 10
D8202 N8202 0 diode
R8203 N8202 N8203 10
D8203 N8203 0 diode
R8204 N8203 N8204 10
D8204 N8204 0 diode
R8205 N8204 N8205 10
D8205 N8205 0 diode
R8206 N8205 N8206 10
D8206 N8206 0 diode
R8207 N8206 N8207 10
D8207 N8207 0 diode
R8208 N8207 N8208 10
D8208 N8208 0 diode
R8209 N8208 N8209 10
D8209 N8209 0 diode
R8210 N8209 N8210 10
D8210 N8210 0 diode
R8211 N8210 N8211 10
D8211 N8211 0 diode
R8212 N8211 N8212 10
D8212 N8212 0 diode
R8213 N8212 N8213 10
D8213 N8213 0 diode
R8214 N8213 N8214 10
D8214 N8214 0 diode
R8215 N8214 N8215 10
D8215 N8215 0 diode
R8216 N8215 N8216 10
D8216 N8216 0 diode
R8217 N8216 N8217 10
D8217 N8217 0 diode
R8218 N8217 N8218 10
D8218 N8218 0 diode
R8219 N8218 N8219 10
D8219 N8219 0 diode
R8220 N8219 N8220 10
D8220 N8220 0 diode
R8221 N8220 N8221 10
D8221 N8221 0 diode
R8222 N8221 N8222 10
D8222 N8222 0 diode
R8223 N8222 N8223 10
D8223 N8223 0 diode
R8224 N8223 N8224 10
D8224 N8224 0 diode
R8225 N8224 N8225 10
D8225 N8225 0 diode
R8226 N8225 N8226 10
D8226 N8226 0 diode
R8227 N8226 N8227 10
D8227 N8227 0 diode
R8228 N8227 N8228 10
D8228 N8228 0 diode
R8229 N8228 N8229 10
D8229 N8229 0 diode
R8230 N8229 N8230 10
D8230 N8230 0 diode
R8231 N8230 N8231 10
D8231 N8231 0 diode
R8232 N8231 N8232 10
D8232 N8232 0 diode
R8233 N8232 N8233 10
D8233 N8233 0 diode
R8234 N8233 N8234 10
D8234 N8234 0 diode
R8235 N8234 N8235 10
D8235 N8235 0 diode
R8236 N8235 N8236 10
D8236 N8236 0 diode
R8237 N8236 N8237 10
D8237 N8237 0 diode
R8238 N8237 N8238 10
D8238 N8238 0 diode
R8239 N8238 N8239 10
D8239 N8239 0 diode
R8240 N8239 N8240 10
D8240 N8240 0 diode
R8241 N8240 N8241 10
D8241 N8241 0 diode
R8242 N8241 N8242 10
D8242 N8242 0 diode
R8243 N8242 N8243 10
D8243 N8243 0 diode
R8244 N8243 N8244 10
D8244 N8244 0 diode
R8245 N8244 N8245 10
D8245 N8245 0 diode
R8246 N8245 N8246 10
D8246 N8246 0 diode
R8247 N8246 N8247 10
D8247 N8247 0 diode
R8248 N8247 N8248 10
D8248 N8248 0 diode
R8249 N8248 N8249 10
D8249 N8249 0 diode
R8250 N8249 N8250 10
D8250 N8250 0 diode
R8251 N8250 N8251 10
D8251 N8251 0 diode
R8252 N8251 N8252 10
D8252 N8252 0 diode
R8253 N8252 N8253 10
D8253 N8253 0 diode
R8254 N8253 N8254 10
D8254 N8254 0 diode
R8255 N8254 N8255 10
D8255 N8255 0 diode
R8256 N8255 N8256 10
D8256 N8256 0 diode
R8257 N8256 N8257 10
D8257 N8257 0 diode
R8258 N8257 N8258 10
D8258 N8258 0 diode
R8259 N8258 N8259 10
D8259 N8259 0 diode
R8260 N8259 N8260 10
D8260 N8260 0 diode
R8261 N8260 N8261 10
D8261 N8261 0 diode
R8262 N8261 N8262 10
D8262 N8262 0 diode
R8263 N8262 N8263 10
D8263 N8263 0 diode
R8264 N8263 N8264 10
D8264 N8264 0 diode
R8265 N8264 N8265 10
D8265 N8265 0 diode
R8266 N8265 N8266 10
D8266 N8266 0 diode
R8267 N8266 N8267 10
D8267 N8267 0 diode
R8268 N8267 N8268 10
D8268 N8268 0 diode
R8269 N8268 N8269 10
D8269 N8269 0 diode
R8270 N8269 N8270 10
D8270 N8270 0 diode
R8271 N8270 N8271 10
D8271 N8271 0 diode
R8272 N8271 N8272 10
D8272 N8272 0 diode
R8273 N8272 N8273 10
D8273 N8273 0 diode
R8274 N8273 N8274 10
D8274 N8274 0 diode
R8275 N8274 N8275 10
D8275 N8275 0 diode
R8276 N8275 N8276 10
D8276 N8276 0 diode
R8277 N8276 N8277 10
D8277 N8277 0 diode
R8278 N8277 N8278 10
D8278 N8278 0 diode
R8279 N8278 N8279 10
D8279 N8279 0 diode
R8280 N8279 N8280 10
D8280 N8280 0 diode
R8281 N8280 N8281 10
D8281 N8281 0 diode
R8282 N8281 N8282 10
D8282 N8282 0 diode
R8283 N8282 N8283 10
D8283 N8283 0 diode
R8284 N8283 N8284 10
D8284 N8284 0 diode
R8285 N8284 N8285 10
D8285 N8285 0 diode
R8286 N8285 N8286 10
D8286 N8286 0 diode
R8287 N8286 N8287 10
D8287 N8287 0 diode
R8288 N8287 N8288 10
D8288 N8288 0 diode
R8289 N8288 N8289 10
D8289 N8289 0 diode
R8290 N8289 N8290 10
D8290 N8290 0 diode
R8291 N8290 N8291 10
D8291 N8291 0 diode
R8292 N8291 N8292 10
D8292 N8292 0 diode
R8293 N8292 N8293 10
D8293 N8293 0 diode
R8294 N8293 N8294 10
D8294 N8294 0 diode
R8295 N8294 N8295 10
D8295 N8295 0 diode
R8296 N8295 N8296 10
D8296 N8296 0 diode
R8297 N8296 N8297 10
D8297 N8297 0 diode
R8298 N8297 N8298 10
D8298 N8298 0 diode
R8299 N8298 N8299 10
D8299 N8299 0 diode
R8300 N8299 N8300 10
D8300 N8300 0 diode
R8301 N8300 N8301 10
D8301 N8301 0 diode
R8302 N8301 N8302 10
D8302 N8302 0 diode
R8303 N8302 N8303 10
D8303 N8303 0 diode
R8304 N8303 N8304 10
D8304 N8304 0 diode
R8305 N8304 N8305 10
D8305 N8305 0 diode
R8306 N8305 N8306 10
D8306 N8306 0 diode
R8307 N8306 N8307 10
D8307 N8307 0 diode
R8308 N8307 N8308 10
D8308 N8308 0 diode
R8309 N8308 N8309 10
D8309 N8309 0 diode
R8310 N8309 N8310 10
D8310 N8310 0 diode
R8311 N8310 N8311 10
D8311 N8311 0 diode
R8312 N8311 N8312 10
D8312 N8312 0 diode
R8313 N8312 N8313 10
D8313 N8313 0 diode
R8314 N8313 N8314 10
D8314 N8314 0 diode
R8315 N8314 N8315 10
D8315 N8315 0 diode
R8316 N8315 N8316 10
D8316 N8316 0 diode
R8317 N8316 N8317 10
D8317 N8317 0 diode
R8318 N8317 N8318 10
D8318 N8318 0 diode
R8319 N8318 N8319 10
D8319 N8319 0 diode
R8320 N8319 N8320 10
D8320 N8320 0 diode
R8321 N8320 N8321 10
D8321 N8321 0 diode
R8322 N8321 N8322 10
D8322 N8322 0 diode
R8323 N8322 N8323 10
D8323 N8323 0 diode
R8324 N8323 N8324 10
D8324 N8324 0 diode
R8325 N8324 N8325 10
D8325 N8325 0 diode
R8326 N8325 N8326 10
D8326 N8326 0 diode
R8327 N8326 N8327 10
D8327 N8327 0 diode
R8328 N8327 N8328 10
D8328 N8328 0 diode
R8329 N8328 N8329 10
D8329 N8329 0 diode
R8330 N8329 N8330 10
D8330 N8330 0 diode
R8331 N8330 N8331 10
D8331 N8331 0 diode
R8332 N8331 N8332 10
D8332 N8332 0 diode
R8333 N8332 N8333 10
D8333 N8333 0 diode
R8334 N8333 N8334 10
D8334 N8334 0 diode
R8335 N8334 N8335 10
D8335 N8335 0 diode
R8336 N8335 N8336 10
D8336 N8336 0 diode
R8337 N8336 N8337 10
D8337 N8337 0 diode
R8338 N8337 N8338 10
D8338 N8338 0 diode
R8339 N8338 N8339 10
D8339 N8339 0 diode
R8340 N8339 N8340 10
D8340 N8340 0 diode
R8341 N8340 N8341 10
D8341 N8341 0 diode
R8342 N8341 N8342 10
D8342 N8342 0 diode
R8343 N8342 N8343 10
D8343 N8343 0 diode
R8344 N8343 N8344 10
D8344 N8344 0 diode
R8345 N8344 N8345 10
D8345 N8345 0 diode
R8346 N8345 N8346 10
D8346 N8346 0 diode
R8347 N8346 N8347 10
D8347 N8347 0 diode
R8348 N8347 N8348 10
D8348 N8348 0 diode
R8349 N8348 N8349 10
D8349 N8349 0 diode
R8350 N8349 N8350 10
D8350 N8350 0 diode
R8351 N8350 N8351 10
D8351 N8351 0 diode
R8352 N8351 N8352 10
D8352 N8352 0 diode
R8353 N8352 N8353 10
D8353 N8353 0 diode
R8354 N8353 N8354 10
D8354 N8354 0 diode
R8355 N8354 N8355 10
D8355 N8355 0 diode
R8356 N8355 N8356 10
D8356 N8356 0 diode
R8357 N8356 N8357 10
D8357 N8357 0 diode
R8358 N8357 N8358 10
D8358 N8358 0 diode
R8359 N8358 N8359 10
D8359 N8359 0 diode
R8360 N8359 N8360 10
D8360 N8360 0 diode
R8361 N8360 N8361 10
D8361 N8361 0 diode
R8362 N8361 N8362 10
D8362 N8362 0 diode
R8363 N8362 N8363 10
D8363 N8363 0 diode
R8364 N8363 N8364 10
D8364 N8364 0 diode
R8365 N8364 N8365 10
D8365 N8365 0 diode
R8366 N8365 N8366 10
D8366 N8366 0 diode
R8367 N8366 N8367 10
D8367 N8367 0 diode
R8368 N8367 N8368 10
D8368 N8368 0 diode
R8369 N8368 N8369 10
D8369 N8369 0 diode
R8370 N8369 N8370 10
D8370 N8370 0 diode
R8371 N8370 N8371 10
D8371 N8371 0 diode
R8372 N8371 N8372 10
D8372 N8372 0 diode
R8373 N8372 N8373 10
D8373 N8373 0 diode
R8374 N8373 N8374 10
D8374 N8374 0 diode
R8375 N8374 N8375 10
D8375 N8375 0 diode
R8376 N8375 N8376 10
D8376 N8376 0 diode
R8377 N8376 N8377 10
D8377 N8377 0 diode
R8378 N8377 N8378 10
D8378 N8378 0 diode
R8379 N8378 N8379 10
D8379 N8379 0 diode
R8380 N8379 N8380 10
D8380 N8380 0 diode
R8381 N8380 N8381 10
D8381 N8381 0 diode
R8382 N8381 N8382 10
D8382 N8382 0 diode
R8383 N8382 N8383 10
D8383 N8383 0 diode
R8384 N8383 N8384 10
D8384 N8384 0 diode
R8385 N8384 N8385 10
D8385 N8385 0 diode
R8386 N8385 N8386 10
D8386 N8386 0 diode
R8387 N8386 N8387 10
D8387 N8387 0 diode
R8388 N8387 N8388 10
D8388 N8388 0 diode
R8389 N8388 N8389 10
D8389 N8389 0 diode
R8390 N8389 N8390 10
D8390 N8390 0 diode
R8391 N8390 N8391 10
D8391 N8391 0 diode
R8392 N8391 N8392 10
D8392 N8392 0 diode
R8393 N8392 N8393 10
D8393 N8393 0 diode
R8394 N8393 N8394 10
D8394 N8394 0 diode
R8395 N8394 N8395 10
D8395 N8395 0 diode
R8396 N8395 N8396 10
D8396 N8396 0 diode
R8397 N8396 N8397 10
D8397 N8397 0 diode
R8398 N8397 N8398 10
D8398 N8398 0 diode
R8399 N8398 N8399 10
D8399 N8399 0 diode
R8400 N8399 N8400 10
D8400 N8400 0 diode
R8401 N8400 N8401 10
D8401 N8401 0 diode
R8402 N8401 N8402 10
D8402 N8402 0 diode
R8403 N8402 N8403 10
D8403 N8403 0 diode
R8404 N8403 N8404 10
D8404 N8404 0 diode
R8405 N8404 N8405 10
D8405 N8405 0 diode
R8406 N8405 N8406 10
D8406 N8406 0 diode
R8407 N8406 N8407 10
D8407 N8407 0 diode
R8408 N8407 N8408 10
D8408 N8408 0 diode
R8409 N8408 N8409 10
D8409 N8409 0 diode
R8410 N8409 N8410 10
D8410 N8410 0 diode
R8411 N8410 N8411 10
D8411 N8411 0 diode
R8412 N8411 N8412 10
D8412 N8412 0 diode
R8413 N8412 N8413 10
D8413 N8413 0 diode
R8414 N8413 N8414 10
D8414 N8414 0 diode
R8415 N8414 N8415 10
D8415 N8415 0 diode
R8416 N8415 N8416 10
D8416 N8416 0 diode
R8417 N8416 N8417 10
D8417 N8417 0 diode
R8418 N8417 N8418 10
D8418 N8418 0 diode
R8419 N8418 N8419 10
D8419 N8419 0 diode
R8420 N8419 N8420 10
D8420 N8420 0 diode
R8421 N8420 N8421 10
D8421 N8421 0 diode
R8422 N8421 N8422 10
D8422 N8422 0 diode
R8423 N8422 N8423 10
D8423 N8423 0 diode
R8424 N8423 N8424 10
D8424 N8424 0 diode
R8425 N8424 N8425 10
D8425 N8425 0 diode
R8426 N8425 N8426 10
D8426 N8426 0 diode
R8427 N8426 N8427 10
D8427 N8427 0 diode
R8428 N8427 N8428 10
D8428 N8428 0 diode
R8429 N8428 N8429 10
D8429 N8429 0 diode
R8430 N8429 N8430 10
D8430 N8430 0 diode
R8431 N8430 N8431 10
D8431 N8431 0 diode
R8432 N8431 N8432 10
D8432 N8432 0 diode
R8433 N8432 N8433 10
D8433 N8433 0 diode
R8434 N8433 N8434 10
D8434 N8434 0 diode
R8435 N8434 N8435 10
D8435 N8435 0 diode
R8436 N8435 N8436 10
D8436 N8436 0 diode
R8437 N8436 N8437 10
D8437 N8437 0 diode
R8438 N8437 N8438 10
D8438 N8438 0 diode
R8439 N8438 N8439 10
D8439 N8439 0 diode
R8440 N8439 N8440 10
D8440 N8440 0 diode
R8441 N8440 N8441 10
D8441 N8441 0 diode
R8442 N8441 N8442 10
D8442 N8442 0 diode
R8443 N8442 N8443 10
D8443 N8443 0 diode
R8444 N8443 N8444 10
D8444 N8444 0 diode
R8445 N8444 N8445 10
D8445 N8445 0 diode
R8446 N8445 N8446 10
D8446 N8446 0 diode
R8447 N8446 N8447 10
D8447 N8447 0 diode
R8448 N8447 N8448 10
D8448 N8448 0 diode
R8449 N8448 N8449 10
D8449 N8449 0 diode
R8450 N8449 N8450 10
D8450 N8450 0 diode
R8451 N8450 N8451 10
D8451 N8451 0 diode
R8452 N8451 N8452 10
D8452 N8452 0 diode
R8453 N8452 N8453 10
D8453 N8453 0 diode
R8454 N8453 N8454 10
D8454 N8454 0 diode
R8455 N8454 N8455 10
D8455 N8455 0 diode
R8456 N8455 N8456 10
D8456 N8456 0 diode
R8457 N8456 N8457 10
D8457 N8457 0 diode
R8458 N8457 N8458 10
D8458 N8458 0 diode
R8459 N8458 N8459 10
D8459 N8459 0 diode
R8460 N8459 N8460 10
D8460 N8460 0 diode
R8461 N8460 N8461 10
D8461 N8461 0 diode
R8462 N8461 N8462 10
D8462 N8462 0 diode
R8463 N8462 N8463 10
D8463 N8463 0 diode
R8464 N8463 N8464 10
D8464 N8464 0 diode
R8465 N8464 N8465 10
D8465 N8465 0 diode
R8466 N8465 N8466 10
D8466 N8466 0 diode
R8467 N8466 N8467 10
D8467 N8467 0 diode
R8468 N8467 N8468 10
D8468 N8468 0 diode
R8469 N8468 N8469 10
D8469 N8469 0 diode
R8470 N8469 N8470 10
D8470 N8470 0 diode
R8471 N8470 N8471 10
D8471 N8471 0 diode
R8472 N8471 N8472 10
D8472 N8472 0 diode
R8473 N8472 N8473 10
D8473 N8473 0 diode
R8474 N8473 N8474 10
D8474 N8474 0 diode
R8475 N8474 N8475 10
D8475 N8475 0 diode
R8476 N8475 N8476 10
D8476 N8476 0 diode
R8477 N8476 N8477 10
D8477 N8477 0 diode
R8478 N8477 N8478 10
D8478 N8478 0 diode
R8479 N8478 N8479 10
D8479 N8479 0 diode
R8480 N8479 N8480 10
D8480 N8480 0 diode
R8481 N8480 N8481 10
D8481 N8481 0 diode
R8482 N8481 N8482 10
D8482 N8482 0 diode
R8483 N8482 N8483 10
D8483 N8483 0 diode
R8484 N8483 N8484 10
D8484 N8484 0 diode
R8485 N8484 N8485 10
D8485 N8485 0 diode
R8486 N8485 N8486 10
D8486 N8486 0 diode
R8487 N8486 N8487 10
D8487 N8487 0 diode
R8488 N8487 N8488 10
D8488 N8488 0 diode
R8489 N8488 N8489 10
D8489 N8489 0 diode
R8490 N8489 N8490 10
D8490 N8490 0 diode
R8491 N8490 N8491 10
D8491 N8491 0 diode
R8492 N8491 N8492 10
D8492 N8492 0 diode
R8493 N8492 N8493 10
D8493 N8493 0 diode
R8494 N8493 N8494 10
D8494 N8494 0 diode
R8495 N8494 N8495 10
D8495 N8495 0 diode
R8496 N8495 N8496 10
D8496 N8496 0 diode
R8497 N8496 N8497 10
D8497 N8497 0 diode
R8498 N8497 N8498 10
D8498 N8498 0 diode
R8499 N8498 N8499 10
D8499 N8499 0 diode
R8500 N8499 N8500 10
D8500 N8500 0 diode
R8501 N8500 N8501 10
D8501 N8501 0 diode
R8502 N8501 N8502 10
D8502 N8502 0 diode
R8503 N8502 N8503 10
D8503 N8503 0 diode
R8504 N8503 N8504 10
D8504 N8504 0 diode
R8505 N8504 N8505 10
D8505 N8505 0 diode
R8506 N8505 N8506 10
D8506 N8506 0 diode
R8507 N8506 N8507 10
D8507 N8507 0 diode
R8508 N8507 N8508 10
D8508 N8508 0 diode
R8509 N8508 N8509 10
D8509 N8509 0 diode
R8510 N8509 N8510 10
D8510 N8510 0 diode
R8511 N8510 N8511 10
D8511 N8511 0 diode
R8512 N8511 N8512 10
D8512 N8512 0 diode
R8513 N8512 N8513 10
D8513 N8513 0 diode
R8514 N8513 N8514 10
D8514 N8514 0 diode
R8515 N8514 N8515 10
D8515 N8515 0 diode
R8516 N8515 N8516 10
D8516 N8516 0 diode
R8517 N8516 N8517 10
D8517 N8517 0 diode
R8518 N8517 N8518 10
D8518 N8518 0 diode
R8519 N8518 N8519 10
D8519 N8519 0 diode
R8520 N8519 N8520 10
D8520 N8520 0 diode
R8521 N8520 N8521 10
D8521 N8521 0 diode
R8522 N8521 N8522 10
D8522 N8522 0 diode
R8523 N8522 N8523 10
D8523 N8523 0 diode
R8524 N8523 N8524 10
D8524 N8524 0 diode
R8525 N8524 N8525 10
D8525 N8525 0 diode
R8526 N8525 N8526 10
D8526 N8526 0 diode
R8527 N8526 N8527 10
D8527 N8527 0 diode
R8528 N8527 N8528 10
D8528 N8528 0 diode
R8529 N8528 N8529 10
D8529 N8529 0 diode
R8530 N8529 N8530 10
D8530 N8530 0 diode
R8531 N8530 N8531 10
D8531 N8531 0 diode
R8532 N8531 N8532 10
D8532 N8532 0 diode
R8533 N8532 N8533 10
D8533 N8533 0 diode
R8534 N8533 N8534 10
D8534 N8534 0 diode
R8535 N8534 N8535 10
D8535 N8535 0 diode
R8536 N8535 N8536 10
D8536 N8536 0 diode
R8537 N8536 N8537 10
D8537 N8537 0 diode
R8538 N8537 N8538 10
D8538 N8538 0 diode
R8539 N8538 N8539 10
D8539 N8539 0 diode
R8540 N8539 N8540 10
D8540 N8540 0 diode
R8541 N8540 N8541 10
D8541 N8541 0 diode
R8542 N8541 N8542 10
D8542 N8542 0 diode
R8543 N8542 N8543 10
D8543 N8543 0 diode
R8544 N8543 N8544 10
D8544 N8544 0 diode
R8545 N8544 N8545 10
D8545 N8545 0 diode
R8546 N8545 N8546 10
D8546 N8546 0 diode
R8547 N8546 N8547 10
D8547 N8547 0 diode
R8548 N8547 N8548 10
D8548 N8548 0 diode
R8549 N8548 N8549 10
D8549 N8549 0 diode
R8550 N8549 N8550 10
D8550 N8550 0 diode
R8551 N8550 N8551 10
D8551 N8551 0 diode
R8552 N8551 N8552 10
D8552 N8552 0 diode
R8553 N8552 N8553 10
D8553 N8553 0 diode
R8554 N8553 N8554 10
D8554 N8554 0 diode
R8555 N8554 N8555 10
D8555 N8555 0 diode
R8556 N8555 N8556 10
D8556 N8556 0 diode
R8557 N8556 N8557 10
D8557 N8557 0 diode
R8558 N8557 N8558 10
D8558 N8558 0 diode
R8559 N8558 N8559 10
D8559 N8559 0 diode
R8560 N8559 N8560 10
D8560 N8560 0 diode
R8561 N8560 N8561 10
D8561 N8561 0 diode
R8562 N8561 N8562 10
D8562 N8562 0 diode
R8563 N8562 N8563 10
D8563 N8563 0 diode
R8564 N8563 N8564 10
D8564 N8564 0 diode
R8565 N8564 N8565 10
D8565 N8565 0 diode
R8566 N8565 N8566 10
D8566 N8566 0 diode
R8567 N8566 N8567 10
D8567 N8567 0 diode
R8568 N8567 N8568 10
D8568 N8568 0 diode
R8569 N8568 N8569 10
D8569 N8569 0 diode
R8570 N8569 N8570 10
D8570 N8570 0 diode
R8571 N8570 N8571 10
D8571 N8571 0 diode
R8572 N8571 N8572 10
D8572 N8572 0 diode
R8573 N8572 N8573 10
D8573 N8573 0 diode
R8574 N8573 N8574 10
D8574 N8574 0 diode
R8575 N8574 N8575 10
D8575 N8575 0 diode
R8576 N8575 N8576 10
D8576 N8576 0 diode
R8577 N8576 N8577 10
D8577 N8577 0 diode
R8578 N8577 N8578 10
D8578 N8578 0 diode
R8579 N8578 N8579 10
D8579 N8579 0 diode
R8580 N8579 N8580 10
D8580 N8580 0 diode
R8581 N8580 N8581 10
D8581 N8581 0 diode
R8582 N8581 N8582 10
D8582 N8582 0 diode
R8583 N8582 N8583 10
D8583 N8583 0 diode
R8584 N8583 N8584 10
D8584 N8584 0 diode
R8585 N8584 N8585 10
D8585 N8585 0 diode
R8586 N8585 N8586 10
D8586 N8586 0 diode
R8587 N8586 N8587 10
D8587 N8587 0 diode
R8588 N8587 N8588 10
D8588 N8588 0 diode
R8589 N8588 N8589 10
D8589 N8589 0 diode
R8590 N8589 N8590 10
D8590 N8590 0 diode
R8591 N8590 N8591 10
D8591 N8591 0 diode
R8592 N8591 N8592 10
D8592 N8592 0 diode
R8593 N8592 N8593 10
D8593 N8593 0 diode
R8594 N8593 N8594 10
D8594 N8594 0 diode
R8595 N8594 N8595 10
D8595 N8595 0 diode
R8596 N8595 N8596 10
D8596 N8596 0 diode
R8597 N8596 N8597 10
D8597 N8597 0 diode
R8598 N8597 N8598 10
D8598 N8598 0 diode
R8599 N8598 N8599 10
D8599 N8599 0 diode
R8600 N8599 N8600 10
D8600 N8600 0 diode
R8601 N8600 N8601 10
D8601 N8601 0 diode
R8602 N8601 N8602 10
D8602 N8602 0 diode
R8603 N8602 N8603 10
D8603 N8603 0 diode
R8604 N8603 N8604 10
D8604 N8604 0 diode
R8605 N8604 N8605 10
D8605 N8605 0 diode
R8606 N8605 N8606 10
D8606 N8606 0 diode
R8607 N8606 N8607 10
D8607 N8607 0 diode
R8608 N8607 N8608 10
D8608 N8608 0 diode
R8609 N8608 N8609 10
D8609 N8609 0 diode
R8610 N8609 N8610 10
D8610 N8610 0 diode
R8611 N8610 N8611 10
D8611 N8611 0 diode
R8612 N8611 N8612 10
D8612 N8612 0 diode
R8613 N8612 N8613 10
D8613 N8613 0 diode
R8614 N8613 N8614 10
D8614 N8614 0 diode
R8615 N8614 N8615 10
D8615 N8615 0 diode
R8616 N8615 N8616 10
D8616 N8616 0 diode
R8617 N8616 N8617 10
D8617 N8617 0 diode
R8618 N8617 N8618 10
D8618 N8618 0 diode
R8619 N8618 N8619 10
D8619 N8619 0 diode
R8620 N8619 N8620 10
D8620 N8620 0 diode
R8621 N8620 N8621 10
D8621 N8621 0 diode
R8622 N8621 N8622 10
D8622 N8622 0 diode
R8623 N8622 N8623 10
D8623 N8623 0 diode
R8624 N8623 N8624 10
D8624 N8624 0 diode
R8625 N8624 N8625 10
D8625 N8625 0 diode
R8626 N8625 N8626 10
D8626 N8626 0 diode
R8627 N8626 N8627 10
D8627 N8627 0 diode
R8628 N8627 N8628 10
D8628 N8628 0 diode
R8629 N8628 N8629 10
D8629 N8629 0 diode
R8630 N8629 N8630 10
D8630 N8630 0 diode
R8631 N8630 N8631 10
D8631 N8631 0 diode
R8632 N8631 N8632 10
D8632 N8632 0 diode
R8633 N8632 N8633 10
D8633 N8633 0 diode
R8634 N8633 N8634 10
D8634 N8634 0 diode
R8635 N8634 N8635 10
D8635 N8635 0 diode
R8636 N8635 N8636 10
D8636 N8636 0 diode
R8637 N8636 N8637 10
D8637 N8637 0 diode
R8638 N8637 N8638 10
D8638 N8638 0 diode
R8639 N8638 N8639 10
D8639 N8639 0 diode
R8640 N8639 N8640 10
D8640 N8640 0 diode
R8641 N8640 N8641 10
D8641 N8641 0 diode
R8642 N8641 N8642 10
D8642 N8642 0 diode
R8643 N8642 N8643 10
D8643 N8643 0 diode
R8644 N8643 N8644 10
D8644 N8644 0 diode
R8645 N8644 N8645 10
D8645 N8645 0 diode
R8646 N8645 N8646 10
D8646 N8646 0 diode
R8647 N8646 N8647 10
D8647 N8647 0 diode
R8648 N8647 N8648 10
D8648 N8648 0 diode
R8649 N8648 N8649 10
D8649 N8649 0 diode
R8650 N8649 N8650 10
D8650 N8650 0 diode
R8651 N8650 N8651 10
D8651 N8651 0 diode
R8652 N8651 N8652 10
D8652 N8652 0 diode
R8653 N8652 N8653 10
D8653 N8653 0 diode
R8654 N8653 N8654 10
D8654 N8654 0 diode
R8655 N8654 N8655 10
D8655 N8655 0 diode
R8656 N8655 N8656 10
D8656 N8656 0 diode
R8657 N8656 N8657 10
D8657 N8657 0 diode
R8658 N8657 N8658 10
D8658 N8658 0 diode
R8659 N8658 N8659 10
D8659 N8659 0 diode
R8660 N8659 N8660 10
D8660 N8660 0 diode
R8661 N8660 N8661 10
D8661 N8661 0 diode
R8662 N8661 N8662 10
D8662 N8662 0 diode
R8663 N8662 N8663 10
D8663 N8663 0 diode
R8664 N8663 N8664 10
D8664 N8664 0 diode
R8665 N8664 N8665 10
D8665 N8665 0 diode
R8666 N8665 N8666 10
D8666 N8666 0 diode
R8667 N8666 N8667 10
D8667 N8667 0 diode
R8668 N8667 N8668 10
D8668 N8668 0 diode
R8669 N8668 N8669 10
D8669 N8669 0 diode
R8670 N8669 N8670 10
D8670 N8670 0 diode
R8671 N8670 N8671 10
D8671 N8671 0 diode
R8672 N8671 N8672 10
D8672 N8672 0 diode
R8673 N8672 N8673 10
D8673 N8673 0 diode
R8674 N8673 N8674 10
D8674 N8674 0 diode
R8675 N8674 N8675 10
D8675 N8675 0 diode
R8676 N8675 N8676 10
D8676 N8676 0 diode
R8677 N8676 N8677 10
D8677 N8677 0 diode
R8678 N8677 N8678 10
D8678 N8678 0 diode
R8679 N8678 N8679 10
D8679 N8679 0 diode
R8680 N8679 N8680 10
D8680 N8680 0 diode
R8681 N8680 N8681 10
D8681 N8681 0 diode
R8682 N8681 N8682 10
D8682 N8682 0 diode
R8683 N8682 N8683 10
D8683 N8683 0 diode
R8684 N8683 N8684 10
D8684 N8684 0 diode
R8685 N8684 N8685 10
D8685 N8685 0 diode
R8686 N8685 N8686 10
D8686 N8686 0 diode
R8687 N8686 N8687 10
D8687 N8687 0 diode
R8688 N8687 N8688 10
D8688 N8688 0 diode
R8689 N8688 N8689 10
D8689 N8689 0 diode
R8690 N8689 N8690 10
D8690 N8690 0 diode
R8691 N8690 N8691 10
D8691 N8691 0 diode
R8692 N8691 N8692 10
D8692 N8692 0 diode
R8693 N8692 N8693 10
D8693 N8693 0 diode
R8694 N8693 N8694 10
D8694 N8694 0 diode
R8695 N8694 N8695 10
D8695 N8695 0 diode
R8696 N8695 N8696 10
D8696 N8696 0 diode
R8697 N8696 N8697 10
D8697 N8697 0 diode
R8698 N8697 N8698 10
D8698 N8698 0 diode
R8699 N8698 N8699 10
D8699 N8699 0 diode
R8700 N8699 N8700 10
D8700 N8700 0 diode
R8701 N8700 N8701 10
D8701 N8701 0 diode
R8702 N8701 N8702 10
D8702 N8702 0 diode
R8703 N8702 N8703 10
D8703 N8703 0 diode
R8704 N8703 N8704 10
D8704 N8704 0 diode
R8705 N8704 N8705 10
D8705 N8705 0 diode
R8706 N8705 N8706 10
D8706 N8706 0 diode
R8707 N8706 N8707 10
D8707 N8707 0 diode
R8708 N8707 N8708 10
D8708 N8708 0 diode
R8709 N8708 N8709 10
D8709 N8709 0 diode
R8710 N8709 N8710 10
D8710 N8710 0 diode
R8711 N8710 N8711 10
D8711 N8711 0 diode
R8712 N8711 N8712 10
D8712 N8712 0 diode
R8713 N8712 N8713 10
D8713 N8713 0 diode
R8714 N8713 N8714 10
D8714 N8714 0 diode
R8715 N8714 N8715 10
D8715 N8715 0 diode
R8716 N8715 N8716 10
D8716 N8716 0 diode
R8717 N8716 N8717 10
D8717 N8717 0 diode
R8718 N8717 N8718 10
D8718 N8718 0 diode
R8719 N8718 N8719 10
D8719 N8719 0 diode
R8720 N8719 N8720 10
D8720 N8720 0 diode
R8721 N8720 N8721 10
D8721 N8721 0 diode
R8722 N8721 N8722 10
D8722 N8722 0 diode
R8723 N8722 N8723 10
D8723 N8723 0 diode
R8724 N8723 N8724 10
D8724 N8724 0 diode
R8725 N8724 N8725 10
D8725 N8725 0 diode
R8726 N8725 N8726 10
D8726 N8726 0 diode
R8727 N8726 N8727 10
D8727 N8727 0 diode
R8728 N8727 N8728 10
D8728 N8728 0 diode
R8729 N8728 N8729 10
D8729 N8729 0 diode
R8730 N8729 N8730 10
D8730 N8730 0 diode
R8731 N8730 N8731 10
D8731 N8731 0 diode
R8732 N8731 N8732 10
D8732 N8732 0 diode
R8733 N8732 N8733 10
D8733 N8733 0 diode
R8734 N8733 N8734 10
D8734 N8734 0 diode
R8735 N8734 N8735 10
D8735 N8735 0 diode
R8736 N8735 N8736 10
D8736 N8736 0 diode
R8737 N8736 N8737 10
D8737 N8737 0 diode
R8738 N8737 N8738 10
D8738 N8738 0 diode
R8739 N8738 N8739 10
D8739 N8739 0 diode
R8740 N8739 N8740 10
D8740 N8740 0 diode
R8741 N8740 N8741 10
D8741 N8741 0 diode
R8742 N8741 N8742 10
D8742 N8742 0 diode
R8743 N8742 N8743 10
D8743 N8743 0 diode
R8744 N8743 N8744 10
D8744 N8744 0 diode
R8745 N8744 N8745 10
D8745 N8745 0 diode
R8746 N8745 N8746 10
D8746 N8746 0 diode
R8747 N8746 N8747 10
D8747 N8747 0 diode
R8748 N8747 N8748 10
D8748 N8748 0 diode
R8749 N8748 N8749 10
D8749 N8749 0 diode
R8750 N8749 N8750 10
D8750 N8750 0 diode
R8751 N8750 N8751 10
D8751 N8751 0 diode
R8752 N8751 N8752 10
D8752 N8752 0 diode
R8753 N8752 N8753 10
D8753 N8753 0 diode
R8754 N8753 N8754 10
D8754 N8754 0 diode
R8755 N8754 N8755 10
D8755 N8755 0 diode
R8756 N8755 N8756 10
D8756 N8756 0 diode
R8757 N8756 N8757 10
D8757 N8757 0 diode
R8758 N8757 N8758 10
D8758 N8758 0 diode
R8759 N8758 N8759 10
D8759 N8759 0 diode
R8760 N8759 N8760 10
D8760 N8760 0 diode
R8761 N8760 N8761 10
D8761 N8761 0 diode
R8762 N8761 N8762 10
D8762 N8762 0 diode
R8763 N8762 N8763 10
D8763 N8763 0 diode
R8764 N8763 N8764 10
D8764 N8764 0 diode
R8765 N8764 N8765 10
D8765 N8765 0 diode
R8766 N8765 N8766 10
D8766 N8766 0 diode
R8767 N8766 N8767 10
D8767 N8767 0 diode
R8768 N8767 N8768 10
D8768 N8768 0 diode
R8769 N8768 N8769 10
D8769 N8769 0 diode
R8770 N8769 N8770 10
D8770 N8770 0 diode
R8771 N8770 N8771 10
D8771 N8771 0 diode
R8772 N8771 N8772 10
D8772 N8772 0 diode
R8773 N8772 N8773 10
D8773 N8773 0 diode
R8774 N8773 N8774 10
D8774 N8774 0 diode
R8775 N8774 N8775 10
D8775 N8775 0 diode
R8776 N8775 N8776 10
D8776 N8776 0 diode
R8777 N8776 N8777 10
D8777 N8777 0 diode
R8778 N8777 N8778 10
D8778 N8778 0 diode
R8779 N8778 N8779 10
D8779 N8779 0 diode
R8780 N8779 N8780 10
D8780 N8780 0 diode
R8781 N8780 N8781 10
D8781 N8781 0 diode
R8782 N8781 N8782 10
D8782 N8782 0 diode
R8783 N8782 N8783 10
D8783 N8783 0 diode
R8784 N8783 N8784 10
D8784 N8784 0 diode
R8785 N8784 N8785 10
D8785 N8785 0 diode
R8786 N8785 N8786 10
D8786 N8786 0 diode
R8787 N8786 N8787 10
D8787 N8787 0 diode
R8788 N8787 N8788 10
D8788 N8788 0 diode
R8789 N8788 N8789 10
D8789 N8789 0 diode
R8790 N8789 N8790 10
D8790 N8790 0 diode
R8791 N8790 N8791 10
D8791 N8791 0 diode
R8792 N8791 N8792 10
D8792 N8792 0 diode
R8793 N8792 N8793 10
D8793 N8793 0 diode
R8794 N8793 N8794 10
D8794 N8794 0 diode
R8795 N8794 N8795 10
D8795 N8795 0 diode
R8796 N8795 N8796 10
D8796 N8796 0 diode
R8797 N8796 N8797 10
D8797 N8797 0 diode
R8798 N8797 N8798 10
D8798 N8798 0 diode
R8799 N8798 N8799 10
D8799 N8799 0 diode
R8800 N8799 N8800 10
D8800 N8800 0 diode
R8801 N8800 N8801 10
D8801 N8801 0 diode
R8802 N8801 N8802 10
D8802 N8802 0 diode
R8803 N8802 N8803 10
D8803 N8803 0 diode
R8804 N8803 N8804 10
D8804 N8804 0 diode
R8805 N8804 N8805 10
D8805 N8805 0 diode
R8806 N8805 N8806 10
D8806 N8806 0 diode
R8807 N8806 N8807 10
D8807 N8807 0 diode
R8808 N8807 N8808 10
D8808 N8808 0 diode
R8809 N8808 N8809 10
D8809 N8809 0 diode
R8810 N8809 N8810 10
D8810 N8810 0 diode
R8811 N8810 N8811 10
D8811 N8811 0 diode
R8812 N8811 N8812 10
D8812 N8812 0 diode
R8813 N8812 N8813 10
D8813 N8813 0 diode
R8814 N8813 N8814 10
D8814 N8814 0 diode
R8815 N8814 N8815 10
D8815 N8815 0 diode
R8816 N8815 N8816 10
D8816 N8816 0 diode
R8817 N8816 N8817 10
D8817 N8817 0 diode
R8818 N8817 N8818 10
D8818 N8818 0 diode
R8819 N8818 N8819 10
D8819 N8819 0 diode
R8820 N8819 N8820 10
D8820 N8820 0 diode
R8821 N8820 N8821 10
D8821 N8821 0 diode
R8822 N8821 N8822 10
D8822 N8822 0 diode
R8823 N8822 N8823 10
D8823 N8823 0 diode
R8824 N8823 N8824 10
D8824 N8824 0 diode
R8825 N8824 N8825 10
D8825 N8825 0 diode
R8826 N8825 N8826 10
D8826 N8826 0 diode
R8827 N8826 N8827 10
D8827 N8827 0 diode
R8828 N8827 N8828 10
D8828 N8828 0 diode
R8829 N8828 N8829 10
D8829 N8829 0 diode
R8830 N8829 N8830 10
D8830 N8830 0 diode
R8831 N8830 N8831 10
D8831 N8831 0 diode
R8832 N8831 N8832 10
D8832 N8832 0 diode
R8833 N8832 N8833 10
D8833 N8833 0 diode
R8834 N8833 N8834 10
D8834 N8834 0 diode
R8835 N8834 N8835 10
D8835 N8835 0 diode
R8836 N8835 N8836 10
D8836 N8836 0 diode
R8837 N8836 N8837 10
D8837 N8837 0 diode
R8838 N8837 N8838 10
D8838 N8838 0 diode
R8839 N8838 N8839 10
D8839 N8839 0 diode
R8840 N8839 N8840 10
D8840 N8840 0 diode
R8841 N8840 N8841 10
D8841 N8841 0 diode
R8842 N8841 N8842 10
D8842 N8842 0 diode
R8843 N8842 N8843 10
D8843 N8843 0 diode
R8844 N8843 N8844 10
D8844 N8844 0 diode
R8845 N8844 N8845 10
D8845 N8845 0 diode
R8846 N8845 N8846 10
D8846 N8846 0 diode
R8847 N8846 N8847 10
D8847 N8847 0 diode
R8848 N8847 N8848 10
D8848 N8848 0 diode
R8849 N8848 N8849 10
D8849 N8849 0 diode
R8850 N8849 N8850 10
D8850 N8850 0 diode
R8851 N8850 N8851 10
D8851 N8851 0 diode
R8852 N8851 N8852 10
D8852 N8852 0 diode
R8853 N8852 N8853 10
D8853 N8853 0 diode
R8854 N8853 N8854 10
D8854 N8854 0 diode
R8855 N8854 N8855 10
D8855 N8855 0 diode
R8856 N8855 N8856 10
D8856 N8856 0 diode
R8857 N8856 N8857 10
D8857 N8857 0 diode
R8858 N8857 N8858 10
D8858 N8858 0 diode
R8859 N8858 N8859 10
D8859 N8859 0 diode
R8860 N8859 N8860 10
D8860 N8860 0 diode
R8861 N8860 N8861 10
D8861 N8861 0 diode
R8862 N8861 N8862 10
D8862 N8862 0 diode
R8863 N8862 N8863 10
D8863 N8863 0 diode
R8864 N8863 N8864 10
D8864 N8864 0 diode
R8865 N8864 N8865 10
D8865 N8865 0 diode
R8866 N8865 N8866 10
D8866 N8866 0 diode
R8867 N8866 N8867 10
D8867 N8867 0 diode
R8868 N8867 N8868 10
D8868 N8868 0 diode
R8869 N8868 N8869 10
D8869 N8869 0 diode
R8870 N8869 N8870 10
D8870 N8870 0 diode
R8871 N8870 N8871 10
D8871 N8871 0 diode
R8872 N8871 N8872 10
D8872 N8872 0 diode
R8873 N8872 N8873 10
D8873 N8873 0 diode
R8874 N8873 N8874 10
D8874 N8874 0 diode
R8875 N8874 N8875 10
D8875 N8875 0 diode
R8876 N8875 N8876 10
D8876 N8876 0 diode
R8877 N8876 N8877 10
D8877 N8877 0 diode
R8878 N8877 N8878 10
D8878 N8878 0 diode
R8879 N8878 N8879 10
D8879 N8879 0 diode
R8880 N8879 N8880 10
D8880 N8880 0 diode
R8881 N8880 N8881 10
D8881 N8881 0 diode
R8882 N8881 N8882 10
D8882 N8882 0 diode
R8883 N8882 N8883 10
D8883 N8883 0 diode
R8884 N8883 N8884 10
D8884 N8884 0 diode
R8885 N8884 N8885 10
D8885 N8885 0 diode
R8886 N8885 N8886 10
D8886 N8886 0 diode
R8887 N8886 N8887 10
D8887 N8887 0 diode
R8888 N8887 N8888 10
D8888 N8888 0 diode
R8889 N8888 N8889 10
D8889 N8889 0 diode
R8890 N8889 N8890 10
D8890 N8890 0 diode
R8891 N8890 N8891 10
D8891 N8891 0 diode
R8892 N8891 N8892 10
D8892 N8892 0 diode
R8893 N8892 N8893 10
D8893 N8893 0 diode
R8894 N8893 N8894 10
D8894 N8894 0 diode
R8895 N8894 N8895 10
D8895 N8895 0 diode
R8896 N8895 N8896 10
D8896 N8896 0 diode
R8897 N8896 N8897 10
D8897 N8897 0 diode
R8898 N8897 N8898 10
D8898 N8898 0 diode
R8899 N8898 N8899 10
D8899 N8899 0 diode
R8900 N8899 N8900 10
D8900 N8900 0 diode
R8901 N8900 N8901 10
D8901 N8901 0 diode
R8902 N8901 N8902 10
D8902 N8902 0 diode
R8903 N8902 N8903 10
D8903 N8903 0 diode
R8904 N8903 N8904 10
D8904 N8904 0 diode
R8905 N8904 N8905 10
D8905 N8905 0 diode
R8906 N8905 N8906 10
D8906 N8906 0 diode
R8907 N8906 N8907 10
D8907 N8907 0 diode
R8908 N8907 N8908 10
D8908 N8908 0 diode
R8909 N8908 N8909 10
D8909 N8909 0 diode
R8910 N8909 N8910 10
D8910 N8910 0 diode
R8911 N8910 N8911 10
D8911 N8911 0 diode
R8912 N8911 N8912 10
D8912 N8912 0 diode
R8913 N8912 N8913 10
D8913 N8913 0 diode
R8914 N8913 N8914 10
D8914 N8914 0 diode
R8915 N8914 N8915 10
D8915 N8915 0 diode
R8916 N8915 N8916 10
D8916 N8916 0 diode
R8917 N8916 N8917 10
D8917 N8917 0 diode
R8918 N8917 N8918 10
D8918 N8918 0 diode
R8919 N8918 N8919 10
D8919 N8919 0 diode
R8920 N8919 N8920 10
D8920 N8920 0 diode
R8921 N8920 N8921 10
D8921 N8921 0 diode
R8922 N8921 N8922 10
D8922 N8922 0 diode
R8923 N8922 N8923 10
D8923 N8923 0 diode
R8924 N8923 N8924 10
D8924 N8924 0 diode
R8925 N8924 N8925 10
D8925 N8925 0 diode
R8926 N8925 N8926 10
D8926 N8926 0 diode
R8927 N8926 N8927 10
D8927 N8927 0 diode
R8928 N8927 N8928 10
D8928 N8928 0 diode
R8929 N8928 N8929 10
D8929 N8929 0 diode
R8930 N8929 N8930 10
D8930 N8930 0 diode
R8931 N8930 N8931 10
D8931 N8931 0 diode
R8932 N8931 N8932 10
D8932 N8932 0 diode
R8933 N8932 N8933 10
D8933 N8933 0 diode
R8934 N8933 N8934 10
D8934 N8934 0 diode
R8935 N8934 N8935 10
D8935 N8935 0 diode
R8936 N8935 N8936 10
D8936 N8936 0 diode
R8937 N8936 N8937 10
D8937 N8937 0 diode
R8938 N8937 N8938 10
D8938 N8938 0 diode
R8939 N8938 N8939 10
D8939 N8939 0 diode
R8940 N8939 N8940 10
D8940 N8940 0 diode
R8941 N8940 N8941 10
D8941 N8941 0 diode
R8942 N8941 N8942 10
D8942 N8942 0 diode
R8943 N8942 N8943 10
D8943 N8943 0 diode
R8944 N8943 N8944 10
D8944 N8944 0 diode
R8945 N8944 N8945 10
D8945 N8945 0 diode
R8946 N8945 N8946 10
D8946 N8946 0 diode
R8947 N8946 N8947 10
D8947 N8947 0 diode
R8948 N8947 N8948 10
D8948 N8948 0 diode
R8949 N8948 N8949 10
D8949 N8949 0 diode
R8950 N8949 N8950 10
D8950 N8950 0 diode
R8951 N8950 N8951 10
D8951 N8951 0 diode
R8952 N8951 N8952 10
D8952 N8952 0 diode
R8953 N8952 N8953 10
D8953 N8953 0 diode
R8954 N8953 N8954 10
D8954 N8954 0 diode
R8955 N8954 N8955 10
D8955 N8955 0 diode
R8956 N8955 N8956 10
D8956 N8956 0 diode
R8957 N8956 N8957 10
D8957 N8957 0 diode
R8958 N8957 N8958 10
D8958 N8958 0 diode
R8959 N8958 N8959 10
D8959 N8959 0 diode
R8960 N8959 N8960 10
D8960 N8960 0 diode
R8961 N8960 N8961 10
D8961 N8961 0 diode
R8962 N8961 N8962 10
D8962 N8962 0 diode
R8963 N8962 N8963 10
D8963 N8963 0 diode
R8964 N8963 N8964 10
D8964 N8964 0 diode
R8965 N8964 N8965 10
D8965 N8965 0 diode
R8966 N8965 N8966 10
D8966 N8966 0 diode
R8967 N8966 N8967 10
D8967 N8967 0 diode
R8968 N8967 N8968 10
D8968 N8968 0 diode
R8969 N8968 N8969 10
D8969 N8969 0 diode
R8970 N8969 N8970 10
D8970 N8970 0 diode
R8971 N8970 N8971 10
D8971 N8971 0 diode
R8972 N8971 N8972 10
D8972 N8972 0 diode
R8973 N8972 N8973 10
D8973 N8973 0 diode
R8974 N8973 N8974 10
D8974 N8974 0 diode
R8975 N8974 N8975 10
D8975 N8975 0 diode
R8976 N8975 N8976 10
D8976 N8976 0 diode
R8977 N8976 N8977 10
D8977 N8977 0 diode
R8978 N8977 N8978 10
D8978 N8978 0 diode
R8979 N8978 N8979 10
D8979 N8979 0 diode
R8980 N8979 N8980 10
D8980 N8980 0 diode
R8981 N8980 N8981 10
D8981 N8981 0 diode
R8982 N8981 N8982 10
D8982 N8982 0 diode
R8983 N8982 N8983 10
D8983 N8983 0 diode
R8984 N8983 N8984 10
D8984 N8984 0 diode
R8985 N8984 N8985 10
D8985 N8985 0 diode
R8986 N8985 N8986 10
D8986 N8986 0 diode
R8987 N8986 N8987 10
D8987 N8987 0 diode
R8988 N8987 N8988 10
D8988 N8988 0 diode
R8989 N8988 N8989 10
D8989 N8989 0 diode
R8990 N8989 N8990 10
D8990 N8990 0 diode
R8991 N8990 N8991 10
D8991 N8991 0 diode
R8992 N8991 N8992 10
D8992 N8992 0 diode
R8993 N8992 N8993 10
D8993 N8993 0 diode
R8994 N8993 N8994 10
D8994 N8994 0 diode
R8995 N8994 N8995 10
D8995 N8995 0 diode
R8996 N8995 N8996 10
D8996 N8996 0 diode
R8997 N8996 N8997 10
D8997 N8997 0 diode
R8998 N8997 N8998 10
D8998 N8998 0 diode
R8999 N8998 N8999 10
D8999 N8999 0 diode
R9000 N8999 N9000 10
D9000 N9000 0 diode
R9001 N9000 N9001 10
D9001 N9001 0 diode
R9002 N9001 N9002 10
D9002 N9002 0 diode
R9003 N9002 N9003 10
D9003 N9003 0 diode
R9004 N9003 N9004 10
D9004 N9004 0 diode
R9005 N9004 N9005 10
D9005 N9005 0 diode
R9006 N9005 N9006 10
D9006 N9006 0 diode
R9007 N9006 N9007 10
D9007 N9007 0 diode
R9008 N9007 N9008 10
D9008 N9008 0 diode
R9009 N9008 N9009 10
D9009 N9009 0 diode
R9010 N9009 N9010 10
D9010 N9010 0 diode
R9011 N9010 N9011 10
D9011 N9011 0 diode
R9012 N9011 N9012 10
D9012 N9012 0 diode
R9013 N9012 N9013 10
D9013 N9013 0 diode
R9014 N9013 N9014 10
D9014 N9014 0 diode
R9015 N9014 N9015 10
D9015 N9015 0 diode
R9016 N9015 N9016 10
D9016 N9016 0 diode
R9017 N9016 N9017 10
D9017 N9017 0 diode
R9018 N9017 N9018 10
D9018 N9018 0 diode
R9019 N9018 N9019 10
D9019 N9019 0 diode
R9020 N9019 N9020 10
D9020 N9020 0 diode
R9021 N9020 N9021 10
D9021 N9021 0 diode
R9022 N9021 N9022 10
D9022 N9022 0 diode
R9023 N9022 N9023 10
D9023 N9023 0 diode
R9024 N9023 N9024 10
D9024 N9024 0 diode
R9025 N9024 N9025 10
D9025 N9025 0 diode
R9026 N9025 N9026 10
D9026 N9026 0 diode
R9027 N9026 N9027 10
D9027 N9027 0 diode
R9028 N9027 N9028 10
D9028 N9028 0 diode
R9029 N9028 N9029 10
D9029 N9029 0 diode
R9030 N9029 N9030 10
D9030 N9030 0 diode
R9031 N9030 N9031 10
D9031 N9031 0 diode
R9032 N9031 N9032 10
D9032 N9032 0 diode
R9033 N9032 N9033 10
D9033 N9033 0 diode
R9034 N9033 N9034 10
D9034 N9034 0 diode
R9035 N9034 N9035 10
D9035 N9035 0 diode
R9036 N9035 N9036 10
D9036 N9036 0 diode
R9037 N9036 N9037 10
D9037 N9037 0 diode
R9038 N9037 N9038 10
D9038 N9038 0 diode
R9039 N9038 N9039 10
D9039 N9039 0 diode
R9040 N9039 N9040 10
D9040 N9040 0 diode
R9041 N9040 N9041 10
D9041 N9041 0 diode
R9042 N9041 N9042 10
D9042 N9042 0 diode
R9043 N9042 N9043 10
D9043 N9043 0 diode
R9044 N9043 N9044 10
D9044 N9044 0 diode
R9045 N9044 N9045 10
D9045 N9045 0 diode
R9046 N9045 N9046 10
D9046 N9046 0 diode
R9047 N9046 N9047 10
D9047 N9047 0 diode
R9048 N9047 N9048 10
D9048 N9048 0 diode
R9049 N9048 N9049 10
D9049 N9049 0 diode
R9050 N9049 N9050 10
D9050 N9050 0 diode
R9051 N9050 N9051 10
D9051 N9051 0 diode
R9052 N9051 N9052 10
D9052 N9052 0 diode
R9053 N9052 N9053 10
D9053 N9053 0 diode
R9054 N9053 N9054 10
D9054 N9054 0 diode
R9055 N9054 N9055 10
D9055 N9055 0 diode
R9056 N9055 N9056 10
D9056 N9056 0 diode
R9057 N9056 N9057 10
D9057 N9057 0 diode
R9058 N9057 N9058 10
D9058 N9058 0 diode
R9059 N9058 N9059 10
D9059 N9059 0 diode
R9060 N9059 N9060 10
D9060 N9060 0 diode
R9061 N9060 N9061 10
D9061 N9061 0 diode
R9062 N9061 N9062 10
D9062 N9062 0 diode
R9063 N9062 N9063 10
D9063 N9063 0 diode
R9064 N9063 N9064 10
D9064 N9064 0 diode
R9065 N9064 N9065 10
D9065 N9065 0 diode
R9066 N9065 N9066 10
D9066 N9066 0 diode
R9067 N9066 N9067 10
D9067 N9067 0 diode
R9068 N9067 N9068 10
D9068 N9068 0 diode
R9069 N9068 N9069 10
D9069 N9069 0 diode
R9070 N9069 N9070 10
D9070 N9070 0 diode
R9071 N9070 N9071 10
D9071 N9071 0 diode
R9072 N9071 N9072 10
D9072 N9072 0 diode
R9073 N9072 N9073 10
D9073 N9073 0 diode
R9074 N9073 N9074 10
D9074 N9074 0 diode
R9075 N9074 N9075 10
D9075 N9075 0 diode
R9076 N9075 N9076 10
D9076 N9076 0 diode
R9077 N9076 N9077 10
D9077 N9077 0 diode
R9078 N9077 N9078 10
D9078 N9078 0 diode
R9079 N9078 N9079 10
D9079 N9079 0 diode
R9080 N9079 N9080 10
D9080 N9080 0 diode
R9081 N9080 N9081 10
D9081 N9081 0 diode
R9082 N9081 N9082 10
D9082 N9082 0 diode
R9083 N9082 N9083 10
D9083 N9083 0 diode
R9084 N9083 N9084 10
D9084 N9084 0 diode
R9085 N9084 N9085 10
D9085 N9085 0 diode
R9086 N9085 N9086 10
D9086 N9086 0 diode
R9087 N9086 N9087 10
D9087 N9087 0 diode
R9088 N9087 N9088 10
D9088 N9088 0 diode
R9089 N9088 N9089 10
D9089 N9089 0 diode
R9090 N9089 N9090 10
D9090 N9090 0 diode
R9091 N9090 N9091 10
D9091 N9091 0 diode
R9092 N9091 N9092 10
D9092 N9092 0 diode
R9093 N9092 N9093 10
D9093 N9093 0 diode
R9094 N9093 N9094 10
D9094 N9094 0 diode
R9095 N9094 N9095 10
D9095 N9095 0 diode
R9096 N9095 N9096 10
D9096 N9096 0 diode
R9097 N9096 N9097 10
D9097 N9097 0 diode
R9098 N9097 N9098 10
D9098 N9098 0 diode
R9099 N9098 N9099 10
D9099 N9099 0 diode
R9100 N9099 N9100 10
D9100 N9100 0 diode
R9101 N9100 N9101 10
D9101 N9101 0 diode
R9102 N9101 N9102 10
D9102 N9102 0 diode
R9103 N9102 N9103 10
D9103 N9103 0 diode
R9104 N9103 N9104 10
D9104 N9104 0 diode
R9105 N9104 N9105 10
D9105 N9105 0 diode
R9106 N9105 N9106 10
D9106 N9106 0 diode
R9107 N9106 N9107 10
D9107 N9107 0 diode
R9108 N9107 N9108 10
D9108 N9108 0 diode
R9109 N9108 N9109 10
D9109 N9109 0 diode
R9110 N9109 N9110 10
D9110 N9110 0 diode
R9111 N9110 N9111 10
D9111 N9111 0 diode
R9112 N9111 N9112 10
D9112 N9112 0 diode
R9113 N9112 N9113 10
D9113 N9113 0 diode
R9114 N9113 N9114 10
D9114 N9114 0 diode
R9115 N9114 N9115 10
D9115 N9115 0 diode
R9116 N9115 N9116 10
D9116 N9116 0 diode
R9117 N9116 N9117 10
D9117 N9117 0 diode
R9118 N9117 N9118 10
D9118 N9118 0 diode
R9119 N9118 N9119 10
D9119 N9119 0 diode
R9120 N9119 N9120 10
D9120 N9120 0 diode
R9121 N9120 N9121 10
D9121 N9121 0 diode
R9122 N9121 N9122 10
D9122 N9122 0 diode
R9123 N9122 N9123 10
D9123 N9123 0 diode
R9124 N9123 N9124 10
D9124 N9124 0 diode
R9125 N9124 N9125 10
D9125 N9125 0 diode
R9126 N9125 N9126 10
D9126 N9126 0 diode
R9127 N9126 N9127 10
D9127 N9127 0 diode
R9128 N9127 N9128 10
D9128 N9128 0 diode
R9129 N9128 N9129 10
D9129 N9129 0 diode
R9130 N9129 N9130 10
D9130 N9130 0 diode
R9131 N9130 N9131 10
D9131 N9131 0 diode
R9132 N9131 N9132 10
D9132 N9132 0 diode
R9133 N9132 N9133 10
D9133 N9133 0 diode
R9134 N9133 N9134 10
D9134 N9134 0 diode
R9135 N9134 N9135 10
D9135 N9135 0 diode
R9136 N9135 N9136 10
D9136 N9136 0 diode
R9137 N9136 N9137 10
D9137 N9137 0 diode
R9138 N9137 N9138 10
D9138 N9138 0 diode
R9139 N9138 N9139 10
D9139 N9139 0 diode
R9140 N9139 N9140 10
D9140 N9140 0 diode
R9141 N9140 N9141 10
D9141 N9141 0 diode
R9142 N9141 N9142 10
D9142 N9142 0 diode
R9143 N9142 N9143 10
D9143 N9143 0 diode
R9144 N9143 N9144 10
D9144 N9144 0 diode
R9145 N9144 N9145 10
D9145 N9145 0 diode
R9146 N9145 N9146 10
D9146 N9146 0 diode
R9147 N9146 N9147 10
D9147 N9147 0 diode
R9148 N9147 N9148 10
D9148 N9148 0 diode
R9149 N9148 N9149 10
D9149 N9149 0 diode
R9150 N9149 N9150 10
D9150 N9150 0 diode
R9151 N9150 N9151 10
D9151 N9151 0 diode
R9152 N9151 N9152 10
D9152 N9152 0 diode
R9153 N9152 N9153 10
D9153 N9153 0 diode
R9154 N9153 N9154 10
D9154 N9154 0 diode
R9155 N9154 N9155 10
D9155 N9155 0 diode
R9156 N9155 N9156 10
D9156 N9156 0 diode
R9157 N9156 N9157 10
D9157 N9157 0 diode
R9158 N9157 N9158 10
D9158 N9158 0 diode
R9159 N9158 N9159 10
D9159 N9159 0 diode
R9160 N9159 N9160 10
D9160 N9160 0 diode
R9161 N9160 N9161 10
D9161 N9161 0 diode
R9162 N9161 N9162 10
D9162 N9162 0 diode
R9163 N9162 N9163 10
D9163 N9163 0 diode
R9164 N9163 N9164 10
D9164 N9164 0 diode
R9165 N9164 N9165 10
D9165 N9165 0 diode
R9166 N9165 N9166 10
D9166 N9166 0 diode
R9167 N9166 N9167 10
D9167 N9167 0 diode
R9168 N9167 N9168 10
D9168 N9168 0 diode
R9169 N9168 N9169 10
D9169 N9169 0 diode
R9170 N9169 N9170 10
D9170 N9170 0 diode
R9171 N9170 N9171 10
D9171 N9171 0 diode
R9172 N9171 N9172 10
D9172 N9172 0 diode
R9173 N9172 N9173 10
D9173 N9173 0 diode
R9174 N9173 N9174 10
D9174 N9174 0 diode
R9175 N9174 N9175 10
D9175 N9175 0 diode
R9176 N9175 N9176 10
D9176 N9176 0 diode
R9177 N9176 N9177 10
D9177 N9177 0 diode
R9178 N9177 N9178 10
D9178 N9178 0 diode
R9179 N9178 N9179 10
D9179 N9179 0 diode
R9180 N9179 N9180 10
D9180 N9180 0 diode
R9181 N9180 N9181 10
D9181 N9181 0 diode
R9182 N9181 N9182 10
D9182 N9182 0 diode
R9183 N9182 N9183 10
D9183 N9183 0 diode
R9184 N9183 N9184 10
D9184 N9184 0 diode
R9185 N9184 N9185 10
D9185 N9185 0 diode
R9186 N9185 N9186 10
D9186 N9186 0 diode
R9187 N9186 N9187 10
D9187 N9187 0 diode
R9188 N9187 N9188 10
D9188 N9188 0 diode
R9189 N9188 N9189 10
D9189 N9189 0 diode
R9190 N9189 N9190 10
D9190 N9190 0 diode
R9191 N9190 N9191 10
D9191 N9191 0 diode
R9192 N9191 N9192 10
D9192 N9192 0 diode
R9193 N9192 N9193 10
D9193 N9193 0 diode
R9194 N9193 N9194 10
D9194 N9194 0 diode
R9195 N9194 N9195 10
D9195 N9195 0 diode
R9196 N9195 N9196 10
D9196 N9196 0 diode
R9197 N9196 N9197 10
D9197 N9197 0 diode
R9198 N9197 N9198 10
D9198 N9198 0 diode
R9199 N9198 N9199 10
D9199 N9199 0 diode
R9200 N9199 N9200 10
D9200 N9200 0 diode
R9201 N9200 N9201 10
D9201 N9201 0 diode
R9202 N9201 N9202 10
D9202 N9202 0 diode
R9203 N9202 N9203 10
D9203 N9203 0 diode
R9204 N9203 N9204 10
D9204 N9204 0 diode
R9205 N9204 N9205 10
D9205 N9205 0 diode
R9206 N9205 N9206 10
D9206 N9206 0 diode
R9207 N9206 N9207 10
D9207 N9207 0 diode
R9208 N9207 N9208 10
D9208 N9208 0 diode
R9209 N9208 N9209 10
D9209 N9209 0 diode
R9210 N9209 N9210 10
D9210 N9210 0 diode
R9211 N9210 N9211 10
D9211 N9211 0 diode
R9212 N9211 N9212 10
D9212 N9212 0 diode
R9213 N9212 N9213 10
D9213 N9213 0 diode
R9214 N9213 N9214 10
D9214 N9214 0 diode
R9215 N9214 N9215 10
D9215 N9215 0 diode
R9216 N9215 N9216 10
D9216 N9216 0 diode
R9217 N9216 N9217 10
D9217 N9217 0 diode
R9218 N9217 N9218 10
D9218 N9218 0 diode
R9219 N9218 N9219 10
D9219 N9219 0 diode
R9220 N9219 N9220 10
D9220 N9220 0 diode
R9221 N9220 N9221 10
D9221 N9221 0 diode
R9222 N9221 N9222 10
D9222 N9222 0 diode
R9223 N9222 N9223 10
D9223 N9223 0 diode
R9224 N9223 N9224 10
D9224 N9224 0 diode
R9225 N9224 N9225 10
D9225 N9225 0 diode
R9226 N9225 N9226 10
D9226 N9226 0 diode
R9227 N9226 N9227 10
D9227 N9227 0 diode
R9228 N9227 N9228 10
D9228 N9228 0 diode
R9229 N9228 N9229 10
D9229 N9229 0 diode
R9230 N9229 N9230 10
D9230 N9230 0 diode
R9231 N9230 N9231 10
D9231 N9231 0 diode
R9232 N9231 N9232 10
D9232 N9232 0 diode
R9233 N9232 N9233 10
D9233 N9233 0 diode
R9234 N9233 N9234 10
D9234 N9234 0 diode
R9235 N9234 N9235 10
D9235 N9235 0 diode
R9236 N9235 N9236 10
D9236 N9236 0 diode
R9237 N9236 N9237 10
D9237 N9237 0 diode
R9238 N9237 N9238 10
D9238 N9238 0 diode
R9239 N9238 N9239 10
D9239 N9239 0 diode
R9240 N9239 N9240 10
D9240 N9240 0 diode
R9241 N9240 N9241 10
D9241 N9241 0 diode
R9242 N9241 N9242 10
D9242 N9242 0 diode
R9243 N9242 N9243 10
D9243 N9243 0 diode
R9244 N9243 N9244 10
D9244 N9244 0 diode
R9245 N9244 N9245 10
D9245 N9245 0 diode
R9246 N9245 N9246 10
D9246 N9246 0 diode
R9247 N9246 N9247 10
D9247 N9247 0 diode
R9248 N9247 N9248 10
D9248 N9248 0 diode
R9249 N9248 N9249 10
D9249 N9249 0 diode
R9250 N9249 N9250 10
D9250 N9250 0 diode
R9251 N9250 N9251 10
D9251 N9251 0 diode
R9252 N9251 N9252 10
D9252 N9252 0 diode
R9253 N9252 N9253 10
D9253 N9253 0 diode
R9254 N9253 N9254 10
D9254 N9254 0 diode
R9255 N9254 N9255 10
D9255 N9255 0 diode
R9256 N9255 N9256 10
D9256 N9256 0 diode
R9257 N9256 N9257 10
D9257 N9257 0 diode
R9258 N9257 N9258 10
D9258 N9258 0 diode
R9259 N9258 N9259 10
D9259 N9259 0 diode
R9260 N9259 N9260 10
D9260 N9260 0 diode
R9261 N9260 N9261 10
D9261 N9261 0 diode
R9262 N9261 N9262 10
D9262 N9262 0 diode
R9263 N9262 N9263 10
D9263 N9263 0 diode
R9264 N9263 N9264 10
D9264 N9264 0 diode
R9265 N9264 N9265 10
D9265 N9265 0 diode
R9266 N9265 N9266 10
D9266 N9266 0 diode
R9267 N9266 N9267 10
D9267 N9267 0 diode
R9268 N9267 N9268 10
D9268 N9268 0 diode
R9269 N9268 N9269 10
D9269 N9269 0 diode
R9270 N9269 N9270 10
D9270 N9270 0 diode
R9271 N9270 N9271 10
D9271 N9271 0 diode
R9272 N9271 N9272 10
D9272 N9272 0 diode
R9273 N9272 N9273 10
D9273 N9273 0 diode
R9274 N9273 N9274 10
D9274 N9274 0 diode
R9275 N9274 N9275 10
D9275 N9275 0 diode
R9276 N9275 N9276 10
D9276 N9276 0 diode
R9277 N9276 N9277 10
D9277 N9277 0 diode
R9278 N9277 N9278 10
D9278 N9278 0 diode
R9279 N9278 N9279 10
D9279 N9279 0 diode
R9280 N9279 N9280 10
D9280 N9280 0 diode
R9281 N9280 N9281 10
D9281 N9281 0 diode
R9282 N9281 N9282 10
D9282 N9282 0 diode
R9283 N9282 N9283 10
D9283 N9283 0 diode
R9284 N9283 N9284 10
D9284 N9284 0 diode
R9285 N9284 N9285 10
D9285 N9285 0 diode
R9286 N9285 N9286 10
D9286 N9286 0 diode
R9287 N9286 N9287 10
D9287 N9287 0 diode
R9288 N9287 N9288 10
D9288 N9288 0 diode
R9289 N9288 N9289 10
D9289 N9289 0 diode
R9290 N9289 N9290 10
D9290 N9290 0 diode
R9291 N9290 N9291 10
D9291 N9291 0 diode
R9292 N9291 N9292 10
D9292 N9292 0 diode
R9293 N9292 N9293 10
D9293 N9293 0 diode
R9294 N9293 N9294 10
D9294 N9294 0 diode
R9295 N9294 N9295 10
D9295 N9295 0 diode
R9296 N9295 N9296 10
D9296 N9296 0 diode
R9297 N9296 N9297 10
D9297 N9297 0 diode
R9298 N9297 N9298 10
D9298 N9298 0 diode
R9299 N9298 N9299 10
D9299 N9299 0 diode
R9300 N9299 N9300 10
D9300 N9300 0 diode
R9301 N9300 N9301 10
D9301 N9301 0 diode
R9302 N9301 N9302 10
D9302 N9302 0 diode
R9303 N9302 N9303 10
D9303 N9303 0 diode
R9304 N9303 N9304 10
D9304 N9304 0 diode
R9305 N9304 N9305 10
D9305 N9305 0 diode
R9306 N9305 N9306 10
D9306 N9306 0 diode
R9307 N9306 N9307 10
D9307 N9307 0 diode
R9308 N9307 N9308 10
D9308 N9308 0 diode
R9309 N9308 N9309 10
D9309 N9309 0 diode
R9310 N9309 N9310 10
D9310 N9310 0 diode
R9311 N9310 N9311 10
D9311 N9311 0 diode
R9312 N9311 N9312 10
D9312 N9312 0 diode
R9313 N9312 N9313 10
D9313 N9313 0 diode
R9314 N9313 N9314 10
D9314 N9314 0 diode
R9315 N9314 N9315 10
D9315 N9315 0 diode
R9316 N9315 N9316 10
D9316 N9316 0 diode
R9317 N9316 N9317 10
D9317 N9317 0 diode
R9318 N9317 N9318 10
D9318 N9318 0 diode
R9319 N9318 N9319 10
D9319 N9319 0 diode
R9320 N9319 N9320 10
D9320 N9320 0 diode
R9321 N9320 N9321 10
D9321 N9321 0 diode
R9322 N9321 N9322 10
D9322 N9322 0 diode
R9323 N9322 N9323 10
D9323 N9323 0 diode
R9324 N9323 N9324 10
D9324 N9324 0 diode
R9325 N9324 N9325 10
D9325 N9325 0 diode
R9326 N9325 N9326 10
D9326 N9326 0 diode
R9327 N9326 N9327 10
D9327 N9327 0 diode
R9328 N9327 N9328 10
D9328 N9328 0 diode
R9329 N9328 N9329 10
D9329 N9329 0 diode
R9330 N9329 N9330 10
D9330 N9330 0 diode
R9331 N9330 N9331 10
D9331 N9331 0 diode
R9332 N9331 N9332 10
D9332 N9332 0 diode
R9333 N9332 N9333 10
D9333 N9333 0 diode
R9334 N9333 N9334 10
D9334 N9334 0 diode
R9335 N9334 N9335 10
D9335 N9335 0 diode
R9336 N9335 N9336 10
D9336 N9336 0 diode
R9337 N9336 N9337 10
D9337 N9337 0 diode
R9338 N9337 N9338 10
D9338 N9338 0 diode
R9339 N9338 N9339 10
D9339 N9339 0 diode
R9340 N9339 N9340 10
D9340 N9340 0 diode
R9341 N9340 N9341 10
D9341 N9341 0 diode
R9342 N9341 N9342 10
D9342 N9342 0 diode
R9343 N9342 N9343 10
D9343 N9343 0 diode
R9344 N9343 N9344 10
D9344 N9344 0 diode
R9345 N9344 N9345 10
D9345 N9345 0 diode
R9346 N9345 N9346 10
D9346 N9346 0 diode
R9347 N9346 N9347 10
D9347 N9347 0 diode
R9348 N9347 N9348 10
D9348 N9348 0 diode
R9349 N9348 N9349 10
D9349 N9349 0 diode
R9350 N9349 N9350 10
D9350 N9350 0 diode
R9351 N9350 N9351 10
D9351 N9351 0 diode
R9352 N9351 N9352 10
D9352 N9352 0 diode
R9353 N9352 N9353 10
D9353 N9353 0 diode
R9354 N9353 N9354 10
D9354 N9354 0 diode
R9355 N9354 N9355 10
D9355 N9355 0 diode
R9356 N9355 N9356 10
D9356 N9356 0 diode
R9357 N9356 N9357 10
D9357 N9357 0 diode
R9358 N9357 N9358 10
D9358 N9358 0 diode
R9359 N9358 N9359 10
D9359 N9359 0 diode
R9360 N9359 N9360 10
D9360 N9360 0 diode
R9361 N9360 N9361 10
D9361 N9361 0 diode
R9362 N9361 N9362 10
D9362 N9362 0 diode
R9363 N9362 N9363 10
D9363 N9363 0 diode
R9364 N9363 N9364 10
D9364 N9364 0 diode
R9365 N9364 N9365 10
D9365 N9365 0 diode
R9366 N9365 N9366 10
D9366 N9366 0 diode
R9367 N9366 N9367 10
D9367 N9367 0 diode
R9368 N9367 N9368 10
D9368 N9368 0 diode
R9369 N9368 N9369 10
D9369 N9369 0 diode
R9370 N9369 N9370 10
D9370 N9370 0 diode
R9371 N9370 N9371 10
D9371 N9371 0 diode
R9372 N9371 N9372 10
D9372 N9372 0 diode
R9373 N9372 N9373 10
D9373 N9373 0 diode
R9374 N9373 N9374 10
D9374 N9374 0 diode
R9375 N9374 N9375 10
D9375 N9375 0 diode
R9376 N9375 N9376 10
D9376 N9376 0 diode
R9377 N9376 N9377 10
D9377 N9377 0 diode
R9378 N9377 N9378 10
D9378 N9378 0 diode
R9379 N9378 N9379 10
D9379 N9379 0 diode
R9380 N9379 N9380 10
D9380 N9380 0 diode
R9381 N9380 N9381 10
D9381 N9381 0 diode
R9382 N9381 N9382 10
D9382 N9382 0 diode
R9383 N9382 N9383 10
D9383 N9383 0 diode
R9384 N9383 N9384 10
D9384 N9384 0 diode
R9385 N9384 N9385 10
D9385 N9385 0 diode
R9386 N9385 N9386 10
D9386 N9386 0 diode
R9387 N9386 N9387 10
D9387 N9387 0 diode
R9388 N9387 N9388 10
D9388 N9388 0 diode
R9389 N9388 N9389 10
D9389 N9389 0 diode
R9390 N9389 N9390 10
D9390 N9390 0 diode
R9391 N9390 N9391 10
D9391 N9391 0 diode
R9392 N9391 N9392 10
D9392 N9392 0 diode
R9393 N9392 N9393 10
D9393 N9393 0 diode
R9394 N9393 N9394 10
D9394 N9394 0 diode
R9395 N9394 N9395 10
D9395 N9395 0 diode
R9396 N9395 N9396 10
D9396 N9396 0 diode
R9397 N9396 N9397 10
D9397 N9397 0 diode
R9398 N9397 N9398 10
D9398 N9398 0 diode
R9399 N9398 N9399 10
D9399 N9399 0 diode
R9400 N9399 N9400 10
D9400 N9400 0 diode
R9401 N9400 N9401 10
D9401 N9401 0 diode
R9402 N9401 N9402 10
D9402 N9402 0 diode
R9403 N9402 N9403 10
D9403 N9403 0 diode
R9404 N9403 N9404 10
D9404 N9404 0 diode
R9405 N9404 N9405 10
D9405 N9405 0 diode
R9406 N9405 N9406 10
D9406 N9406 0 diode
R9407 N9406 N9407 10
D9407 N9407 0 diode
R9408 N9407 N9408 10
D9408 N9408 0 diode
R9409 N9408 N9409 10
D9409 N9409 0 diode
R9410 N9409 N9410 10
D9410 N9410 0 diode
R9411 N9410 N9411 10
D9411 N9411 0 diode
R9412 N9411 N9412 10
D9412 N9412 0 diode
R9413 N9412 N9413 10
D9413 N9413 0 diode
R9414 N9413 N9414 10
D9414 N9414 0 diode
R9415 N9414 N9415 10
D9415 N9415 0 diode
R9416 N9415 N9416 10
D9416 N9416 0 diode
R9417 N9416 N9417 10
D9417 N9417 0 diode
R9418 N9417 N9418 10
D9418 N9418 0 diode
R9419 N9418 N9419 10
D9419 N9419 0 diode
R9420 N9419 N9420 10
D9420 N9420 0 diode
R9421 N9420 N9421 10
D9421 N9421 0 diode
R9422 N9421 N9422 10
D9422 N9422 0 diode
R9423 N9422 N9423 10
D9423 N9423 0 diode
R9424 N9423 N9424 10
D9424 N9424 0 diode
R9425 N9424 N9425 10
D9425 N9425 0 diode
R9426 N9425 N9426 10
D9426 N9426 0 diode
R9427 N9426 N9427 10
D9427 N9427 0 diode
R9428 N9427 N9428 10
D9428 N9428 0 diode
R9429 N9428 N9429 10
D9429 N9429 0 diode
R9430 N9429 N9430 10
D9430 N9430 0 diode
R9431 N9430 N9431 10
D9431 N9431 0 diode
R9432 N9431 N9432 10
D9432 N9432 0 diode
R9433 N9432 N9433 10
D9433 N9433 0 diode
R9434 N9433 N9434 10
D9434 N9434 0 diode
R9435 N9434 N9435 10
D9435 N9435 0 diode
R9436 N9435 N9436 10
D9436 N9436 0 diode
R9437 N9436 N9437 10
D9437 N9437 0 diode
R9438 N9437 N9438 10
D9438 N9438 0 diode
R9439 N9438 N9439 10
D9439 N9439 0 diode
R9440 N9439 N9440 10
D9440 N9440 0 diode
R9441 N9440 N9441 10
D9441 N9441 0 diode
R9442 N9441 N9442 10
D9442 N9442 0 diode
R9443 N9442 N9443 10
D9443 N9443 0 diode
R9444 N9443 N9444 10
D9444 N9444 0 diode
R9445 N9444 N9445 10
D9445 N9445 0 diode
R9446 N9445 N9446 10
D9446 N9446 0 diode
R9447 N9446 N9447 10
D9447 N9447 0 diode
R9448 N9447 N9448 10
D9448 N9448 0 diode
R9449 N9448 N9449 10
D9449 N9449 0 diode
R9450 N9449 N9450 10
D9450 N9450 0 diode
R9451 N9450 N9451 10
D9451 N9451 0 diode
R9452 N9451 N9452 10
D9452 N9452 0 diode
R9453 N9452 N9453 10
D9453 N9453 0 diode
R9454 N9453 N9454 10
D9454 N9454 0 diode
R9455 N9454 N9455 10
D9455 N9455 0 diode
R9456 N9455 N9456 10
D9456 N9456 0 diode
R9457 N9456 N9457 10
D9457 N9457 0 diode
R9458 N9457 N9458 10
D9458 N9458 0 diode
R9459 N9458 N9459 10
D9459 N9459 0 diode
R9460 N9459 N9460 10
D9460 N9460 0 diode
R9461 N9460 N9461 10
D9461 N9461 0 diode
R9462 N9461 N9462 10
D9462 N9462 0 diode
R9463 N9462 N9463 10
D9463 N9463 0 diode
R9464 N9463 N9464 10
D9464 N9464 0 diode
R9465 N9464 N9465 10
D9465 N9465 0 diode
R9466 N9465 N9466 10
D9466 N9466 0 diode
R9467 N9466 N9467 10
D9467 N9467 0 diode
R9468 N9467 N9468 10
D9468 N9468 0 diode
R9469 N9468 N9469 10
D9469 N9469 0 diode
R9470 N9469 N9470 10
D9470 N9470 0 diode
R9471 N9470 N9471 10
D9471 N9471 0 diode
R9472 N9471 N9472 10
D9472 N9472 0 diode
R9473 N9472 N9473 10
D9473 N9473 0 diode
R9474 N9473 N9474 10
D9474 N9474 0 diode
R9475 N9474 N9475 10
D9475 N9475 0 diode
R9476 N9475 N9476 10
D9476 N9476 0 diode
R9477 N9476 N9477 10
D9477 N9477 0 diode
R9478 N9477 N9478 10
D9478 N9478 0 diode
R9479 N9478 N9479 10
D9479 N9479 0 diode
R9480 N9479 N9480 10
D9480 N9480 0 diode
R9481 N9480 N9481 10
D9481 N9481 0 diode
R9482 N9481 N9482 10
D9482 N9482 0 diode
R9483 N9482 N9483 10
D9483 N9483 0 diode
R9484 N9483 N9484 10
D9484 N9484 0 diode
R9485 N9484 N9485 10
D9485 N9485 0 diode
R9486 N9485 N9486 10
D9486 N9486 0 diode
R9487 N9486 N9487 10
D9487 N9487 0 diode
R9488 N9487 N9488 10
D9488 N9488 0 diode
R9489 N9488 N9489 10
D9489 N9489 0 diode
R9490 N9489 N9490 10
D9490 N9490 0 diode
R9491 N9490 N9491 10
D9491 N9491 0 diode
R9492 N9491 N9492 10
D9492 N9492 0 diode
R9493 N9492 N9493 10
D9493 N9493 0 diode
R9494 N9493 N9494 10
D9494 N9494 0 diode
R9495 N9494 N9495 10
D9495 N9495 0 diode
R9496 N9495 N9496 10
D9496 N9496 0 diode
R9497 N9496 N9497 10
D9497 N9497 0 diode
R9498 N9497 N9498 10
D9498 N9498 0 diode
R9499 N9498 N9499 10
D9499 N9499 0 diode
R9500 N9499 N9500 10
D9500 N9500 0 diode
R9501 N9500 N9501 10
D9501 N9501 0 diode
R9502 N9501 N9502 10
D9502 N9502 0 diode
R9503 N9502 N9503 10
D9503 N9503 0 diode
R9504 N9503 N9504 10
D9504 N9504 0 diode
R9505 N9504 N9505 10
D9505 N9505 0 diode
R9506 N9505 N9506 10
D9506 N9506 0 diode
R9507 N9506 N9507 10
D9507 N9507 0 diode
R9508 N9507 N9508 10
D9508 N9508 0 diode
R9509 N9508 N9509 10
D9509 N9509 0 diode
R9510 N9509 N9510 10
D9510 N9510 0 diode
R9511 N9510 N9511 10
D9511 N9511 0 diode
R9512 N9511 N9512 10
D9512 N9512 0 diode
R9513 N9512 N9513 10
D9513 N9513 0 diode
R9514 N9513 N9514 10
D9514 N9514 0 diode
R9515 N9514 N9515 10
D9515 N9515 0 diode
R9516 N9515 N9516 10
D9516 N9516 0 diode
R9517 N9516 N9517 10
D9517 N9517 0 diode
R9518 N9517 N9518 10
D9518 N9518 0 diode
R9519 N9518 N9519 10
D9519 N9519 0 diode
R9520 N9519 N9520 10
D9520 N9520 0 diode
R9521 N9520 N9521 10
D9521 N9521 0 diode
R9522 N9521 N9522 10
D9522 N9522 0 diode
R9523 N9522 N9523 10
D9523 N9523 0 diode
R9524 N9523 N9524 10
D9524 N9524 0 diode
R9525 N9524 N9525 10
D9525 N9525 0 diode
R9526 N9525 N9526 10
D9526 N9526 0 diode
R9527 N9526 N9527 10
D9527 N9527 0 diode
R9528 N9527 N9528 10
D9528 N9528 0 diode
R9529 N9528 N9529 10
D9529 N9529 0 diode
R9530 N9529 N9530 10
D9530 N9530 0 diode
R9531 N9530 N9531 10
D9531 N9531 0 diode
R9532 N9531 N9532 10
D9532 N9532 0 diode
R9533 N9532 N9533 10
D9533 N9533 0 diode
R9534 N9533 N9534 10
D9534 N9534 0 diode
R9535 N9534 N9535 10
D9535 N9535 0 diode
R9536 N9535 N9536 10
D9536 N9536 0 diode
R9537 N9536 N9537 10
D9537 N9537 0 diode
R9538 N9537 N9538 10
D9538 N9538 0 diode
R9539 N9538 N9539 10
D9539 N9539 0 diode
R9540 N9539 N9540 10
D9540 N9540 0 diode
R9541 N9540 N9541 10
D9541 N9541 0 diode
R9542 N9541 N9542 10
D9542 N9542 0 diode
R9543 N9542 N9543 10
D9543 N9543 0 diode
R9544 N9543 N9544 10
D9544 N9544 0 diode
R9545 N9544 N9545 10
D9545 N9545 0 diode
R9546 N9545 N9546 10
D9546 N9546 0 diode
R9547 N9546 N9547 10
D9547 N9547 0 diode
R9548 N9547 N9548 10
D9548 N9548 0 diode
R9549 N9548 N9549 10
D9549 N9549 0 diode
R9550 N9549 N9550 10
D9550 N9550 0 diode
R9551 N9550 N9551 10
D9551 N9551 0 diode
R9552 N9551 N9552 10
D9552 N9552 0 diode
R9553 N9552 N9553 10
D9553 N9553 0 diode
R9554 N9553 N9554 10
D9554 N9554 0 diode
R9555 N9554 N9555 10
D9555 N9555 0 diode
R9556 N9555 N9556 10
D9556 N9556 0 diode
R9557 N9556 N9557 10
D9557 N9557 0 diode
R9558 N9557 N9558 10
D9558 N9558 0 diode
R9559 N9558 N9559 10
D9559 N9559 0 diode
R9560 N9559 N9560 10
D9560 N9560 0 diode
R9561 N9560 N9561 10
D9561 N9561 0 diode
R9562 N9561 N9562 10
D9562 N9562 0 diode
R9563 N9562 N9563 10
D9563 N9563 0 diode
R9564 N9563 N9564 10
D9564 N9564 0 diode
R9565 N9564 N9565 10
D9565 N9565 0 diode
R9566 N9565 N9566 10
D9566 N9566 0 diode
R9567 N9566 N9567 10
D9567 N9567 0 diode
R9568 N9567 N9568 10
D9568 N9568 0 diode
R9569 N9568 N9569 10
D9569 N9569 0 diode
R9570 N9569 N9570 10
D9570 N9570 0 diode
R9571 N9570 N9571 10
D9571 N9571 0 diode
R9572 N9571 N9572 10
D9572 N9572 0 diode
R9573 N9572 N9573 10
D9573 N9573 0 diode
R9574 N9573 N9574 10
D9574 N9574 0 diode
R9575 N9574 N9575 10
D9575 N9575 0 diode
R9576 N9575 N9576 10
D9576 N9576 0 diode
R9577 N9576 N9577 10
D9577 N9577 0 diode
R9578 N9577 N9578 10
D9578 N9578 0 diode
R9579 N9578 N9579 10
D9579 N9579 0 diode
R9580 N9579 N9580 10
D9580 N9580 0 diode
R9581 N9580 N9581 10
D9581 N9581 0 diode
R9582 N9581 N9582 10
D9582 N9582 0 diode
R9583 N9582 N9583 10
D9583 N9583 0 diode
R9584 N9583 N9584 10
D9584 N9584 0 diode
R9585 N9584 N9585 10
D9585 N9585 0 diode
R9586 N9585 N9586 10
D9586 N9586 0 diode
R9587 N9586 N9587 10
D9587 N9587 0 diode
R9588 N9587 N9588 10
D9588 N9588 0 diode
R9589 N9588 N9589 10
D9589 N9589 0 diode
R9590 N9589 N9590 10
D9590 N9590 0 diode
R9591 N9590 N9591 10
D9591 N9591 0 diode
R9592 N9591 N9592 10
D9592 N9592 0 diode
R9593 N9592 N9593 10
D9593 N9593 0 diode
R9594 N9593 N9594 10
D9594 N9594 0 diode
R9595 N9594 N9595 10
D9595 N9595 0 diode
R9596 N9595 N9596 10
D9596 N9596 0 diode
R9597 N9596 N9597 10
D9597 N9597 0 diode
R9598 N9597 N9598 10
D9598 N9598 0 diode
R9599 N9598 N9599 10
D9599 N9599 0 diode
R9600 N9599 N9600 10
D9600 N9600 0 diode
R9601 N9600 N9601 10
D9601 N9601 0 diode
R9602 N9601 N9602 10
D9602 N9602 0 diode
R9603 N9602 N9603 10
D9603 N9603 0 diode
R9604 N9603 N9604 10
D9604 N9604 0 diode
R9605 N9604 N9605 10
D9605 N9605 0 diode
R9606 N9605 N9606 10
D9606 N9606 0 diode
R9607 N9606 N9607 10
D9607 N9607 0 diode
R9608 N9607 N9608 10
D9608 N9608 0 diode
R9609 N9608 N9609 10
D9609 N9609 0 diode
R9610 N9609 N9610 10
D9610 N9610 0 diode
R9611 N9610 N9611 10
D9611 N9611 0 diode
R9612 N9611 N9612 10
D9612 N9612 0 diode
R9613 N9612 N9613 10
D9613 N9613 0 diode
R9614 N9613 N9614 10
D9614 N9614 0 diode
R9615 N9614 N9615 10
D9615 N9615 0 diode
R9616 N9615 N9616 10
D9616 N9616 0 diode
R9617 N9616 N9617 10
D9617 N9617 0 diode
R9618 N9617 N9618 10
D9618 N9618 0 diode
R9619 N9618 N9619 10
D9619 N9619 0 diode
R9620 N9619 N9620 10
D9620 N9620 0 diode
R9621 N9620 N9621 10
D9621 N9621 0 diode
R9622 N9621 N9622 10
D9622 N9622 0 diode
R9623 N9622 N9623 10
D9623 N9623 0 diode
R9624 N9623 N9624 10
D9624 N9624 0 diode
R9625 N9624 N9625 10
D9625 N9625 0 diode
R9626 N9625 N9626 10
D9626 N9626 0 diode
R9627 N9626 N9627 10
D9627 N9627 0 diode
R9628 N9627 N9628 10
D9628 N9628 0 diode
R9629 N9628 N9629 10
D9629 N9629 0 diode
R9630 N9629 N9630 10
D9630 N9630 0 diode
R9631 N9630 N9631 10
D9631 N9631 0 diode
R9632 N9631 N9632 10
D9632 N9632 0 diode
R9633 N9632 N9633 10
D9633 N9633 0 diode
R9634 N9633 N9634 10
D9634 N9634 0 diode
R9635 N9634 N9635 10
D9635 N9635 0 diode
R9636 N9635 N9636 10
D9636 N9636 0 diode
R9637 N9636 N9637 10
D9637 N9637 0 diode
R9638 N9637 N9638 10
D9638 N9638 0 diode
R9639 N9638 N9639 10
D9639 N9639 0 diode
R9640 N9639 N9640 10
D9640 N9640 0 diode
R9641 N9640 N9641 10
D9641 N9641 0 diode
R9642 N9641 N9642 10
D9642 N9642 0 diode
R9643 N9642 N9643 10
D9643 N9643 0 diode
R9644 N9643 N9644 10
D9644 N9644 0 diode
R9645 N9644 N9645 10
D9645 N9645 0 diode
R9646 N9645 N9646 10
D9646 N9646 0 diode
R9647 N9646 N9647 10
D9647 N9647 0 diode
R9648 N9647 N9648 10
D9648 N9648 0 diode
R9649 N9648 N9649 10
D9649 N9649 0 diode
R9650 N9649 N9650 10
D9650 N9650 0 diode
R9651 N9650 N9651 10
D9651 N9651 0 diode
R9652 N9651 N9652 10
D9652 N9652 0 diode
R9653 N9652 N9653 10
D9653 N9653 0 diode
R9654 N9653 N9654 10
D9654 N9654 0 diode
R9655 N9654 N9655 10
D9655 N9655 0 diode
R9656 N9655 N9656 10
D9656 N9656 0 diode
R9657 N9656 N9657 10
D9657 N9657 0 diode
R9658 N9657 N9658 10
D9658 N9658 0 diode
R9659 N9658 N9659 10
D9659 N9659 0 diode
R9660 N9659 N9660 10
D9660 N9660 0 diode
R9661 N9660 N9661 10
D9661 N9661 0 diode
R9662 N9661 N9662 10
D9662 N9662 0 diode
R9663 N9662 N9663 10
D9663 N9663 0 diode
R9664 N9663 N9664 10
D9664 N9664 0 diode
R9665 N9664 N9665 10
D9665 N9665 0 diode
R9666 N9665 N9666 10
D9666 N9666 0 diode
R9667 N9666 N9667 10
D9667 N9667 0 diode
R9668 N9667 N9668 10
D9668 N9668 0 diode
R9669 N9668 N9669 10
D9669 N9669 0 diode
R9670 N9669 N9670 10
D9670 N9670 0 diode
R9671 N9670 N9671 10
D9671 N9671 0 diode
R9672 N9671 N9672 10
D9672 N9672 0 diode
R9673 N9672 N9673 10
D9673 N9673 0 diode
R9674 N9673 N9674 10
D9674 N9674 0 diode
R9675 N9674 N9675 10
D9675 N9675 0 diode
R9676 N9675 N9676 10
D9676 N9676 0 diode
R9677 N9676 N9677 10
D9677 N9677 0 diode
R9678 N9677 N9678 10
D9678 N9678 0 diode
R9679 N9678 N9679 10
D9679 N9679 0 diode
R9680 N9679 N9680 10
D9680 N9680 0 diode
R9681 N9680 N9681 10
D9681 N9681 0 diode
R9682 N9681 N9682 10
D9682 N9682 0 diode
R9683 N9682 N9683 10
D9683 N9683 0 diode
R9684 N9683 N9684 10
D9684 N9684 0 diode
R9685 N9684 N9685 10
D9685 N9685 0 diode
R9686 N9685 N9686 10
D9686 N9686 0 diode
R9687 N9686 N9687 10
D9687 N9687 0 diode
R9688 N9687 N9688 10
D9688 N9688 0 diode
R9689 N9688 N9689 10
D9689 N9689 0 diode
R9690 N9689 N9690 10
D9690 N9690 0 diode
R9691 N9690 N9691 10
D9691 N9691 0 diode
R9692 N9691 N9692 10
D9692 N9692 0 diode
R9693 N9692 N9693 10
D9693 N9693 0 diode
R9694 N9693 N9694 10
D9694 N9694 0 diode
R9695 N9694 N9695 10
D9695 N9695 0 diode
R9696 N9695 N9696 10
D9696 N9696 0 diode
R9697 N9696 N9697 10
D9697 N9697 0 diode
R9698 N9697 N9698 10
D9698 N9698 0 diode
R9699 N9698 N9699 10
D9699 N9699 0 diode
R9700 N9699 N9700 10
D9700 N9700 0 diode
R9701 N9700 N9701 10
D9701 N9701 0 diode
R9702 N9701 N9702 10
D9702 N9702 0 diode
R9703 N9702 N9703 10
D9703 N9703 0 diode
R9704 N9703 N9704 10
D9704 N9704 0 diode
R9705 N9704 N9705 10
D9705 N9705 0 diode
R9706 N9705 N9706 10
D9706 N9706 0 diode
R9707 N9706 N9707 10
D9707 N9707 0 diode
R9708 N9707 N9708 10
D9708 N9708 0 diode
R9709 N9708 N9709 10
D9709 N9709 0 diode
R9710 N9709 N9710 10
D9710 N9710 0 diode
R9711 N9710 N9711 10
D9711 N9711 0 diode
R9712 N9711 N9712 10
D9712 N9712 0 diode
R9713 N9712 N9713 10
D9713 N9713 0 diode
R9714 N9713 N9714 10
D9714 N9714 0 diode
R9715 N9714 N9715 10
D9715 N9715 0 diode
R9716 N9715 N9716 10
D9716 N9716 0 diode
R9717 N9716 N9717 10
D9717 N9717 0 diode
R9718 N9717 N9718 10
D9718 N9718 0 diode
R9719 N9718 N9719 10
D9719 N9719 0 diode
R9720 N9719 N9720 10
D9720 N9720 0 diode
R9721 N9720 N9721 10
D9721 N9721 0 diode
R9722 N9721 N9722 10
D9722 N9722 0 diode
R9723 N9722 N9723 10
D9723 N9723 0 diode
R9724 N9723 N9724 10
D9724 N9724 0 diode
R9725 N9724 N9725 10
D9725 N9725 0 diode
R9726 N9725 N9726 10
D9726 N9726 0 diode
R9727 N9726 N9727 10
D9727 N9727 0 diode
R9728 N9727 N9728 10
D9728 N9728 0 diode
R9729 N9728 N9729 10
D9729 N9729 0 diode
R9730 N9729 N9730 10
D9730 N9730 0 diode
R9731 N9730 N9731 10
D9731 N9731 0 diode
R9732 N9731 N9732 10
D9732 N9732 0 diode
R9733 N9732 N9733 10
D9733 N9733 0 diode
R9734 N9733 N9734 10
D9734 N9734 0 diode
R9735 N9734 N9735 10
D9735 N9735 0 diode
R9736 N9735 N9736 10
D9736 N9736 0 diode
R9737 N9736 N9737 10
D9737 N9737 0 diode
R9738 N9737 N9738 10
D9738 N9738 0 diode
R9739 N9738 N9739 10
D9739 N9739 0 diode
R9740 N9739 N9740 10
D9740 N9740 0 diode
R9741 N9740 N9741 10
D9741 N9741 0 diode
R9742 N9741 N9742 10
D9742 N9742 0 diode
R9743 N9742 N9743 10
D9743 N9743 0 diode
R9744 N9743 N9744 10
D9744 N9744 0 diode
R9745 N9744 N9745 10
D9745 N9745 0 diode
R9746 N9745 N9746 10
D9746 N9746 0 diode
R9747 N9746 N9747 10
D9747 N9747 0 diode
R9748 N9747 N9748 10
D9748 N9748 0 diode
R9749 N9748 N9749 10
D9749 N9749 0 diode
R9750 N9749 N9750 10
D9750 N9750 0 diode
R9751 N9750 N9751 10
D9751 N9751 0 diode
R9752 N9751 N9752 10
D9752 N9752 0 diode
R9753 N9752 N9753 10
D9753 N9753 0 diode
R9754 N9753 N9754 10
D9754 N9754 0 diode
R9755 N9754 N9755 10
D9755 N9755 0 diode
R9756 N9755 N9756 10
D9756 N9756 0 diode
R9757 N9756 N9757 10
D9757 N9757 0 diode
R9758 N9757 N9758 10
D9758 N9758 0 diode
R9759 N9758 N9759 10
D9759 N9759 0 diode
R9760 N9759 N9760 10
D9760 N9760 0 diode
R9761 N9760 N9761 10
D9761 N9761 0 diode
R9762 N9761 N9762 10
D9762 N9762 0 diode
R9763 N9762 N9763 10
D9763 N9763 0 diode
R9764 N9763 N9764 10
D9764 N9764 0 diode
R9765 N9764 N9765 10
D9765 N9765 0 diode
R9766 N9765 N9766 10
D9766 N9766 0 diode
R9767 N9766 N9767 10
D9767 N9767 0 diode
R9768 N9767 N9768 10
D9768 N9768 0 diode
R9769 N9768 N9769 10
D9769 N9769 0 diode
R9770 N9769 N9770 10
D9770 N9770 0 diode
R9771 N9770 N9771 10
D9771 N9771 0 diode
R9772 N9771 N9772 10
D9772 N9772 0 diode
R9773 N9772 N9773 10
D9773 N9773 0 diode
R9774 N9773 N9774 10
D9774 N9774 0 diode
R9775 N9774 N9775 10
D9775 N9775 0 diode
R9776 N9775 N9776 10
D9776 N9776 0 diode
R9777 N9776 N9777 10
D9777 N9777 0 diode
R9778 N9777 N9778 10
D9778 N9778 0 diode
R9779 N9778 N9779 10
D9779 N9779 0 diode
R9780 N9779 N9780 10
D9780 N9780 0 diode
R9781 N9780 N9781 10
D9781 N9781 0 diode
R9782 N9781 N9782 10
D9782 N9782 0 diode
R9783 N9782 N9783 10
D9783 N9783 0 diode
R9784 N9783 N9784 10
D9784 N9784 0 diode
R9785 N9784 N9785 10
D9785 N9785 0 diode
R9786 N9785 N9786 10
D9786 N9786 0 diode
R9787 N9786 N9787 10
D9787 N9787 0 diode
R9788 N9787 N9788 10
D9788 N9788 0 diode
R9789 N9788 N9789 10
D9789 N9789 0 diode
R9790 N9789 N9790 10
D9790 N9790 0 diode
R9791 N9790 N9791 10
D9791 N9791 0 diode
R9792 N9791 N9792 10
D9792 N9792 0 diode
R9793 N9792 N9793 10
D9793 N9793 0 diode
R9794 N9793 N9794 10
D9794 N9794 0 diode
R9795 N9794 N9795 10
D9795 N9795 0 diode
R9796 N9795 N9796 10
D9796 N9796 0 diode
R9797 N9796 N9797 10
D9797 N9797 0 diode
R9798 N9797 N9798 10
D9798 N9798 0 diode
R9799 N9798 N9799 10
D9799 N9799 0 diode
R9800 N9799 N9800 10
D9800 N9800 0 diode
R9801 N9800 N9801 10
D9801 N9801 0 diode
R9802 N9801 N9802 10
D9802 N9802 0 diode
R9803 N9802 N9803 10
D9803 N9803 0 diode
R9804 N9803 N9804 10
D9804 N9804 0 diode
R9805 N9804 N9805 10
D9805 N9805 0 diode
R9806 N9805 N9806 10
D9806 N9806 0 diode
R9807 N9806 N9807 10
D9807 N9807 0 diode
R9808 N9807 N9808 10
D9808 N9808 0 diode
R9809 N9808 N9809 10
D9809 N9809 0 diode
R9810 N9809 N9810 10
D9810 N9810 0 diode
R9811 N9810 N9811 10
D9811 N9811 0 diode
R9812 N9811 N9812 10
D9812 N9812 0 diode
R9813 N9812 N9813 10
D9813 N9813 0 diode
R9814 N9813 N9814 10
D9814 N9814 0 diode
R9815 N9814 N9815 10
D9815 N9815 0 diode
R9816 N9815 N9816 10
D9816 N9816 0 diode
R9817 N9816 N9817 10
D9817 N9817 0 diode
R9818 N9817 N9818 10
D9818 N9818 0 diode
R9819 N9818 N9819 10
D9819 N9819 0 diode
R9820 N9819 N9820 10
D9820 N9820 0 diode
R9821 N9820 N9821 10
D9821 N9821 0 diode
R9822 N9821 N9822 10
D9822 N9822 0 diode
R9823 N9822 N9823 10
D9823 N9823 0 diode
R9824 N9823 N9824 10
D9824 N9824 0 diode
R9825 N9824 N9825 10
D9825 N9825 0 diode
R9826 N9825 N9826 10
D9826 N9826 0 diode
R9827 N9826 N9827 10
D9827 N9827 0 diode
R9828 N9827 N9828 10
D9828 N9828 0 diode
R9829 N9828 N9829 10
D9829 N9829 0 diode
R9830 N9829 N9830 10
D9830 N9830 0 diode
R9831 N9830 N9831 10
D9831 N9831 0 diode
R9832 N9831 N9832 10
D9832 N9832 0 diode
R9833 N9832 N9833 10
D9833 N9833 0 diode
R9834 N9833 N9834 10
D9834 N9834 0 diode
R9835 N9834 N9835 10
D9835 N9835 0 diode
R9836 N9835 N9836 10
D9836 N9836 0 diode
R9837 N9836 N9837 10
D9837 N9837 0 diode
R9838 N9837 N9838 10
D9838 N9838 0 diode
R9839 N9838 N9839 10
D9839 N9839 0 diode
R9840 N9839 N9840 10
D9840 N9840 0 diode
R9841 N9840 N9841 10
D9841 N9841 0 diode
R9842 N9841 N9842 10
D9842 N9842 0 diode
R9843 N9842 N9843 10
D9843 N9843 0 diode
R9844 N9843 N9844 10
D9844 N9844 0 diode
R9845 N9844 N9845 10
D9845 N9845 0 diode
R9846 N9845 N9846 10
D9846 N9846 0 diode
R9847 N9846 N9847 10
D9847 N9847 0 diode
R9848 N9847 N9848 10
D9848 N9848 0 diode
R9849 N9848 N9849 10
D9849 N9849 0 diode
R9850 N9849 N9850 10
D9850 N9850 0 diode
R9851 N9850 N9851 10
D9851 N9851 0 diode
R9852 N9851 N9852 10
D9852 N9852 0 diode
R9853 N9852 N9853 10
D9853 N9853 0 diode
R9854 N9853 N9854 10
D9854 N9854 0 diode
R9855 N9854 N9855 10
D9855 N9855 0 diode
R9856 N9855 N9856 10
D9856 N9856 0 diode
R9857 N9856 N9857 10
D9857 N9857 0 diode
R9858 N9857 N9858 10
D9858 N9858 0 diode
R9859 N9858 N9859 10
D9859 N9859 0 diode
R9860 N9859 N9860 10
D9860 N9860 0 diode
R9861 N9860 N9861 10
D9861 N9861 0 diode
R9862 N9861 N9862 10
D9862 N9862 0 diode
R9863 N9862 N9863 10
D9863 N9863 0 diode
R9864 N9863 N9864 10
D9864 N9864 0 diode
R9865 N9864 N9865 10
D9865 N9865 0 diode
R9866 N9865 N9866 10
D9866 N9866 0 diode
R9867 N9866 N9867 10
D9867 N9867 0 diode
R9868 N9867 N9868 10
D9868 N9868 0 diode
R9869 N9868 N9869 10
D9869 N9869 0 diode
R9870 N9869 N9870 10
D9870 N9870 0 diode
R9871 N9870 N9871 10
D9871 N9871 0 diode
R9872 N9871 N9872 10
D9872 N9872 0 diode
R9873 N9872 N9873 10
D9873 N9873 0 diode
R9874 N9873 N9874 10
D9874 N9874 0 diode
R9875 N9874 N9875 10
D9875 N9875 0 diode
R9876 N9875 N9876 10
D9876 N9876 0 diode
R9877 N9876 N9877 10
D9877 N9877 0 diode
R9878 N9877 N9878 10
D9878 N9878 0 diode
R9879 N9878 N9879 10
D9879 N9879 0 diode
R9880 N9879 N9880 10
D9880 N9880 0 diode
R9881 N9880 N9881 10
D9881 N9881 0 diode
R9882 N9881 N9882 10
D9882 N9882 0 diode
R9883 N9882 N9883 10
D9883 N9883 0 diode
R9884 N9883 N9884 10
D9884 N9884 0 diode
R9885 N9884 N9885 10
D9885 N9885 0 diode
R9886 N9885 N9886 10
D9886 N9886 0 diode
R9887 N9886 N9887 10
D9887 N9887 0 diode
R9888 N9887 N9888 10
D9888 N9888 0 diode
R9889 N9888 N9889 10
D9889 N9889 0 diode
R9890 N9889 N9890 10
D9890 N9890 0 diode
R9891 N9890 N9891 10
D9891 N9891 0 diode
R9892 N9891 N9892 10
D9892 N9892 0 diode
R9893 N9892 N9893 10
D9893 N9893 0 diode
R9894 N9893 N9894 10
D9894 N9894 0 diode
R9895 N9894 N9895 10
D9895 N9895 0 diode
R9896 N9895 N9896 10
D9896 N9896 0 diode
R9897 N9896 N9897 10
D9897 N9897 0 diode
R9898 N9897 N9898 10
D9898 N9898 0 diode
R9899 N9898 N9899 10
D9899 N9899 0 diode
R9900 N9899 N9900 10
D9900 N9900 0 diode
R9901 N9900 N9901 10
D9901 N9901 0 diode
R9902 N9901 N9902 10
D9902 N9902 0 diode
R9903 N9902 N9903 10
D9903 N9903 0 diode
R9904 N9903 N9904 10
D9904 N9904 0 diode
R9905 N9904 N9905 10
D9905 N9905 0 diode
R9906 N9905 N9906 10
D9906 N9906 0 diode
R9907 N9906 N9907 10
D9907 N9907 0 diode
R9908 N9907 N9908 10
D9908 N9908 0 diode
R9909 N9908 N9909 10
D9909 N9909 0 diode
R9910 N9909 N9910 10
D9910 N9910 0 diode
R9911 N9910 N9911 10
D9911 N9911 0 diode
R9912 N9911 N9912 10
D9912 N9912 0 diode
R9913 N9912 N9913 10
D9913 N9913 0 diode
R9914 N9913 N9914 10
D9914 N9914 0 diode
R9915 N9914 N9915 10
D9915 N9915 0 diode
R9916 N9915 N9916 10
D9916 N9916 0 diode
R9917 N9916 N9917 10
D9917 N9917 0 diode
R9918 N9917 N9918 10
D9918 N9918 0 diode
R9919 N9918 N9919 10
D9919 N9919 0 diode
R9920 N9919 N9920 10
D9920 N9920 0 diode
R9921 N9920 N9921 10
D9921 N9921 0 diode
R9922 N9921 N9922 10
D9922 N9922 0 diode
R9923 N9922 N9923 10
D9923 N9923 0 diode
R9924 N9923 N9924 10
D9924 N9924 0 diode
R9925 N9924 N9925 10
D9925 N9925 0 diode
R9926 N9925 N9926 10
D9926 N9926 0 diode
R9927 N9926 N9927 10
D9927 N9927 0 diode
R9928 N9927 N9928 10
D9928 N9928 0 diode
R9929 N9928 N9929 10
D9929 N9929 0 diode
R9930 N9929 N9930 10
D9930 N9930 0 diode
R9931 N9930 N9931 10
D9931 N9931 0 diode
R9932 N9931 N9932 10
D9932 N9932 0 diode
R9933 N9932 N9933 10
D9933 N9933 0 diode
R9934 N9933 N9934 10
D9934 N9934 0 diode
R9935 N9934 N9935 10
D9935 N9935 0 diode
R9936 N9935 N9936 10
D9936 N9936 0 diode
R9937 N9936 N9937 10
D9937 N9937 0 diode
R9938 N9937 N9938 10
D9938 N9938 0 diode
R9939 N9938 N9939 10
D9939 N9939 0 diode
R9940 N9939 N9940 10
D9940 N9940 0 diode
R9941 N9940 N9941 10
D9941 N9941 0 diode
R9942 N9941 N9942 10
D9942 N9942 0 diode
R9943 N9942 N9943 10
D9943 N9943 0 diode
R9944 N9943 N9944 10
D9944 N9944 0 diode
R9945 N9944 N9945 10
D9945 N9945 0 diode
R9946 N9945 N9946 10
D9946 N9946 0 diode
R9947 N9946 N9947 10
D9947 N9947 0 diode
R9948 N9947 N9948 10
D9948 N9948 0 diode
R9949 N9948 N9949 10
D9949 N9949 0 diode
R9950 N9949 N9950 10
D9950 N9950 0 diode
R9951 N9950 N9951 10
D9951 N9951 0 diode
R9952 N9951 N9952 10
D9952 N9952 0 diode
R9953 N9952 N9953 10
D9953 N9953 0 diode
R9954 N9953 N9954 10
D9954 N9954 0 diode
R9955 N9954 N9955 10
D9955 N9955 0 diode
R9956 N9955 N9956 10
D9956 N9956 0 diode
R9957 N9956 N9957 10
D9957 N9957 0 diode
R9958 N9957 N9958 10
D9958 N9958 0 diode
R9959 N9958 N9959 10
D9959 N9959 0 diode
R9960 N9959 N9960 10
D9960 N9960 0 diode
R9961 N9960 N9961 10
D9961 N9961 0 diode
R9962 N9961 N9962 10
D9962 N9962 0 diode
R9963 N9962 N9963 10
D9963 N9963 0 diode
R9964 N9963 N9964 10
D9964 N9964 0 diode
R9965 N9964 N9965 10
D9965 N9965 0 diode
R9966 N9965 N9966 10
D9966 N9966 0 diode
R9967 N9966 N9967 10
D9967 N9967 0 diode
R9968 N9967 N9968 10
D9968 N9968 0 diode
R9969 N9968 N9969 10
D9969 N9969 0 diode
R9970 N9969 N9970 10
D9970 N9970 0 diode
R9971 N9970 N9971 10
D9971 N9971 0 diode
R9972 N9971 N9972 10
D9972 N9972 0 diode
R9973 N9972 N9973 10
D9973 N9973 0 diode
R9974 N9973 N9974 10
D9974 N9974 0 diode
R9975 N9974 N9975 10
D9975 N9975 0 diode
R9976 N9975 N9976 10
D9976 N9976 0 diode
R9977 N9976 N9977 10
D9977 N9977 0 diode
R9978 N9977 N9978 10
D9978 N9978 0 diode
R9979 N9978 N9979 10
D9979 N9979 0 diode
R9980 N9979 N9980 10
D9980 N9980 0 diode
R9981 N9980 N9981 10
D9981 N9981 0 diode
R9982 N9981 N9982 10
D9982 N9982 0 diode
R9983 N9982 N9983 10
D9983 N9983 0 diode
R9984 N9983 N9984 10
D9984 N9984 0 diode
R9985 N9984 N9985 10
D9985 N9985 0 diode
R9986 N9985 N9986 10
D9986 N9986 0 diode
R9987 N9986 N9987 10
D9987 N9987 0 diode
R9988 N9987 N9988 10
D9988 N9988 0 diode
R9989 N9988 N9989 10
D9989 N9989 0 diode
R9990 N9989 N9990 10
D9990 N9990 0 diode
R9991 N9990 N9991 10
D9991 N9991 0 diode
R9992 N9991 N9992 10
D9992 N9992 0 diode
R9993 N9992 N9993 10
D9993 N9993 0 diode
R9994 N9993 N9994 10
D9994 N9994 0 diode
R9995 N9994 N9995 10
D9995 N9995 0 diode
R9996 N9995 N9996 10
D9996 N9996 0 diode
R9997 N9996 N9997 10
D9997 N9997 0 diode
R9998 N9997 N9998 10
D9998 N9998 0 diode
R9999 N9998 N9999 10
D9999 N9999 0 diode
R10000 N9999 N10000 10
D10000 N10000 0 diode
R10001 N10000 N10001 10
D10001 N10001 0 diode
R10002 N10001 N10002 10
D10002 N10002 0 diode
R10003 N10002 N10003 10
D10003 N10003 0 diode
R10004 N10003 N10004 10
D10004 N10004 0 diode
R10005 N10004 N10005 10
D10005 N10005 0 diode
R10006 N10005 N10006 10
D10006 N10006 0 diode
R10007 N10006 N10007 10
D10007 N10007 0 diode
R10008 N10007 N10008 10
D10008 N10008 0 diode
R10009 N10008 N10009 10
D10009 N10009 0 diode
R10010 N10009 N10010 10
D10010 N10010 0 diode
R10011 N10010 N10011 10
D10011 N10011 0 diode
R10012 N10011 N10012 10
D10012 N10012 0 diode
R10013 N10012 N10013 10
D10013 N10013 0 diode
R10014 N10013 N10014 10
D10014 N10014 0 diode
R10015 N10014 N10015 10
D10015 N10015 0 diode
R10016 N10015 N10016 10
D10016 N10016 0 diode
R10017 N10016 N10017 10
D10017 N10017 0 diode
R10018 N10017 N10018 10
D10018 N10018 0 diode
R10019 N10018 N10019 10
D10019 N10019 0 diode
R10020 N10019 N10020 10
D10020 N10020 0 diode
R10021 N10020 N10021 10
D10021 N10021 0 diode
R10022 N10021 N10022 10
D10022 N10022 0 diode
R10023 N10022 N10023 10
D10023 N10023 0 diode
R10024 N10023 N10024 10
D10024 N10024 0 diode
R10025 N10024 N10025 10
D10025 N10025 0 diode
R10026 N10025 N10026 10
D10026 N10026 0 diode
R10027 N10026 N10027 10
D10027 N10027 0 diode
R10028 N10027 N10028 10
D10028 N10028 0 diode
R10029 N10028 N10029 10
D10029 N10029 0 diode
R10030 N10029 N10030 10
D10030 N10030 0 diode
R10031 N10030 N10031 10
D10031 N10031 0 diode
R10032 N10031 N10032 10
D10032 N10032 0 diode
R10033 N10032 N10033 10
D10033 N10033 0 diode
R10034 N10033 N10034 10
D10034 N10034 0 diode
R10035 N10034 N10035 10
D10035 N10035 0 diode
R10036 N10035 N10036 10
D10036 N10036 0 diode
R10037 N10036 N10037 10
D10037 N10037 0 diode
R10038 N10037 N10038 10
D10038 N10038 0 diode
R10039 N10038 N10039 10
D10039 N10039 0 diode
R10040 N10039 N10040 10
D10040 N10040 0 diode
R10041 N10040 N10041 10
D10041 N10041 0 diode
R10042 N10041 N10042 10
D10042 N10042 0 diode
R10043 N10042 N10043 10
D10043 N10043 0 diode
R10044 N10043 N10044 10
D10044 N10044 0 diode
R10045 N10044 N10045 10
D10045 N10045 0 diode
R10046 N10045 N10046 10
D10046 N10046 0 diode
R10047 N10046 N10047 10
D10047 N10047 0 diode
R10048 N10047 N10048 10
D10048 N10048 0 diode
R10049 N10048 N10049 10
D10049 N10049 0 diode
R10050 N10049 N10050 10
D10050 N10050 0 diode
R10051 N10050 N10051 10
D10051 N10051 0 diode
R10052 N10051 N10052 10
D10052 N10052 0 diode
R10053 N10052 N10053 10
D10053 N10053 0 diode
R10054 N10053 N10054 10
D10054 N10054 0 diode
R10055 N10054 N10055 10
D10055 N10055 0 diode
R10056 N10055 N10056 10
D10056 N10056 0 diode
R10057 N10056 N10057 10
D10057 N10057 0 diode
R10058 N10057 N10058 10
D10058 N10058 0 diode
R10059 N10058 N10059 10
D10059 N10059 0 diode
R10060 N10059 N10060 10
D10060 N10060 0 diode
R10061 N10060 N10061 10
D10061 N10061 0 diode
R10062 N10061 N10062 10
D10062 N10062 0 diode
R10063 N10062 N10063 10
D10063 N10063 0 diode
R10064 N10063 N10064 10
D10064 N10064 0 diode
R10065 N10064 N10065 10
D10065 N10065 0 diode
R10066 N10065 N10066 10
D10066 N10066 0 diode
R10067 N10066 N10067 10
D10067 N10067 0 diode
R10068 N10067 N10068 10
D10068 N10068 0 diode
R10069 N10068 N10069 10
D10069 N10069 0 diode
R10070 N10069 N10070 10
D10070 N10070 0 diode
R10071 N10070 N10071 10
D10071 N10071 0 diode
R10072 N10071 N10072 10
D10072 N10072 0 diode
R10073 N10072 N10073 10
D10073 N10073 0 diode
R10074 N10073 N10074 10
D10074 N10074 0 diode
R10075 N10074 N10075 10
D10075 N10075 0 diode
R10076 N10075 N10076 10
D10076 N10076 0 diode
R10077 N10076 N10077 10
D10077 N10077 0 diode
R10078 N10077 N10078 10
D10078 N10078 0 diode
R10079 N10078 N10079 10
D10079 N10079 0 diode
R10080 N10079 N10080 10
D10080 N10080 0 diode
R10081 N10080 N10081 10
D10081 N10081 0 diode
R10082 N10081 N10082 10
D10082 N10082 0 diode
R10083 N10082 N10083 10
D10083 N10083 0 diode
R10084 N10083 N10084 10
D10084 N10084 0 diode
R10085 N10084 N10085 10
D10085 N10085 0 diode
R10086 N10085 N10086 10
D10086 N10086 0 diode
R10087 N10086 N10087 10
D10087 N10087 0 diode
R10088 N10087 N10088 10
D10088 N10088 0 diode
R10089 N10088 N10089 10
D10089 N10089 0 diode
R10090 N10089 N10090 10
D10090 N10090 0 diode
R10091 N10090 N10091 10
D10091 N10091 0 diode
R10092 N10091 N10092 10
D10092 N10092 0 diode
R10093 N10092 N10093 10
D10093 N10093 0 diode
R10094 N10093 N10094 10
D10094 N10094 0 diode
R10095 N10094 N10095 10
D10095 N10095 0 diode
R10096 N10095 N10096 10
D10096 N10096 0 diode
R10097 N10096 N10097 10
D10097 N10097 0 diode
R10098 N10097 N10098 10
D10098 N10098 0 diode
R10099 N10098 N10099 10
D10099 N10099 0 diode
R10100 N10099 N10100 10
D10100 N10100 0 diode
R10101 N10100 N10101 10
D10101 N10101 0 diode
R10102 N10101 N10102 10
D10102 N10102 0 diode
R10103 N10102 N10103 10
D10103 N10103 0 diode
R10104 N10103 N10104 10
D10104 N10104 0 diode
R10105 N10104 N10105 10
D10105 N10105 0 diode
R10106 N10105 N10106 10
D10106 N10106 0 diode
R10107 N10106 N10107 10
D10107 N10107 0 diode
R10108 N10107 N10108 10
D10108 N10108 0 diode
R10109 N10108 N10109 10
D10109 N10109 0 diode
R10110 N10109 N10110 10
D10110 N10110 0 diode
R10111 N10110 N10111 10
D10111 N10111 0 diode
R10112 N10111 N10112 10
D10112 N10112 0 diode
R10113 N10112 N10113 10
D10113 N10113 0 diode
R10114 N10113 N10114 10
D10114 N10114 0 diode
R10115 N10114 N10115 10
D10115 N10115 0 diode
R10116 N10115 N10116 10
D10116 N10116 0 diode
R10117 N10116 N10117 10
D10117 N10117 0 diode
R10118 N10117 N10118 10
D10118 N10118 0 diode
R10119 N10118 N10119 10
D10119 N10119 0 diode
R10120 N10119 N10120 10
D10120 N10120 0 diode
R10121 N10120 N10121 10
D10121 N10121 0 diode
R10122 N10121 N10122 10
D10122 N10122 0 diode
R10123 N10122 N10123 10
D10123 N10123 0 diode
R10124 N10123 N10124 10
D10124 N10124 0 diode
R10125 N10124 N10125 10
D10125 N10125 0 diode
R10126 N10125 N10126 10
D10126 N10126 0 diode
R10127 N10126 N10127 10
D10127 N10127 0 diode
R10128 N10127 N10128 10
D10128 N10128 0 diode
R10129 N10128 N10129 10
D10129 N10129 0 diode
R10130 N10129 N10130 10
D10130 N10130 0 diode
R10131 N10130 N10131 10
D10131 N10131 0 diode
R10132 N10131 N10132 10
D10132 N10132 0 diode
R10133 N10132 N10133 10
D10133 N10133 0 diode
R10134 N10133 N10134 10
D10134 N10134 0 diode
R10135 N10134 N10135 10
D10135 N10135 0 diode
R10136 N10135 N10136 10
D10136 N10136 0 diode
R10137 N10136 N10137 10
D10137 N10137 0 diode
R10138 N10137 N10138 10
D10138 N10138 0 diode
R10139 N10138 N10139 10
D10139 N10139 0 diode
R10140 N10139 N10140 10
D10140 N10140 0 diode
R10141 N10140 N10141 10
D10141 N10141 0 diode
R10142 N10141 N10142 10
D10142 N10142 0 diode
R10143 N10142 N10143 10
D10143 N10143 0 diode
R10144 N10143 N10144 10
D10144 N10144 0 diode
R10145 N10144 N10145 10
D10145 N10145 0 diode
R10146 N10145 N10146 10
D10146 N10146 0 diode
R10147 N10146 N10147 10
D10147 N10147 0 diode
R10148 N10147 N10148 10
D10148 N10148 0 diode
R10149 N10148 N10149 10
D10149 N10149 0 diode
R10150 N10149 N10150 10
D10150 N10150 0 diode
R10151 N10150 N10151 10
D10151 N10151 0 diode
R10152 N10151 N10152 10
D10152 N10152 0 diode
R10153 N10152 N10153 10
D10153 N10153 0 diode
R10154 N10153 N10154 10
D10154 N10154 0 diode
R10155 N10154 N10155 10
D10155 N10155 0 diode
R10156 N10155 N10156 10
D10156 N10156 0 diode
R10157 N10156 N10157 10
D10157 N10157 0 diode
R10158 N10157 N10158 10
D10158 N10158 0 diode
R10159 N10158 N10159 10
D10159 N10159 0 diode
R10160 N10159 N10160 10
D10160 N10160 0 diode
R10161 N10160 N10161 10
D10161 N10161 0 diode
R10162 N10161 N10162 10
D10162 N10162 0 diode
R10163 N10162 N10163 10
D10163 N10163 0 diode
R10164 N10163 N10164 10
D10164 N10164 0 diode
R10165 N10164 N10165 10
D10165 N10165 0 diode
R10166 N10165 N10166 10
D10166 N10166 0 diode
R10167 N10166 N10167 10
D10167 N10167 0 diode
R10168 N10167 N10168 10
D10168 N10168 0 diode
R10169 N10168 N10169 10
D10169 N10169 0 diode
R10170 N10169 N10170 10
D10170 N10170 0 diode
R10171 N10170 N10171 10
D10171 N10171 0 diode
R10172 N10171 N10172 10
D10172 N10172 0 diode
R10173 N10172 N10173 10
D10173 N10173 0 diode
R10174 N10173 N10174 10
D10174 N10174 0 diode
R10175 N10174 N10175 10
D10175 N10175 0 diode
R10176 N10175 N10176 10
D10176 N10176 0 diode
R10177 N10176 N10177 10
D10177 N10177 0 diode
R10178 N10177 N10178 10
D10178 N10178 0 diode
R10179 N10178 N10179 10
D10179 N10179 0 diode
R10180 N10179 N10180 10
D10180 N10180 0 diode
R10181 N10180 N10181 10
D10181 N10181 0 diode
R10182 N10181 N10182 10
D10182 N10182 0 diode
R10183 N10182 N10183 10
D10183 N10183 0 diode
R10184 N10183 N10184 10
D10184 N10184 0 diode
R10185 N10184 N10185 10
D10185 N10185 0 diode
R10186 N10185 N10186 10
D10186 N10186 0 diode
R10187 N10186 N10187 10
D10187 N10187 0 diode
R10188 N10187 N10188 10
D10188 N10188 0 diode
R10189 N10188 N10189 10
D10189 N10189 0 diode
R10190 N10189 N10190 10
D10190 N10190 0 diode
R10191 N10190 N10191 10
D10191 N10191 0 diode
R10192 N10191 N10192 10
D10192 N10192 0 diode
R10193 N10192 N10193 10
D10193 N10193 0 diode
R10194 N10193 N10194 10
D10194 N10194 0 diode
R10195 N10194 N10195 10
D10195 N10195 0 diode
R10196 N10195 N10196 10
D10196 N10196 0 diode
R10197 N10196 N10197 10
D10197 N10197 0 diode
R10198 N10197 N10198 10
D10198 N10198 0 diode
R10199 N10198 N10199 10
D10199 N10199 0 diode
R10200 N10199 N10200 10
D10200 N10200 0 diode
R10201 N10200 N10201 10
D10201 N10201 0 diode
R10202 N10201 N10202 10
D10202 N10202 0 diode
R10203 N10202 N10203 10
D10203 N10203 0 diode
R10204 N10203 N10204 10
D10204 N10204 0 diode
R10205 N10204 N10205 10
D10205 N10205 0 diode
R10206 N10205 N10206 10
D10206 N10206 0 diode
R10207 N10206 N10207 10
D10207 N10207 0 diode
R10208 N10207 N10208 10
D10208 N10208 0 diode
R10209 N10208 N10209 10
D10209 N10209 0 diode
R10210 N10209 N10210 10
D10210 N10210 0 diode
R10211 N10210 N10211 10
D10211 N10211 0 diode
R10212 N10211 N10212 10
D10212 N10212 0 diode
R10213 N10212 N10213 10
D10213 N10213 0 diode
R10214 N10213 N10214 10
D10214 N10214 0 diode
R10215 N10214 N10215 10
D10215 N10215 0 diode
R10216 N10215 N10216 10
D10216 N10216 0 diode
R10217 N10216 N10217 10
D10217 N10217 0 diode
R10218 N10217 N10218 10
D10218 N10218 0 diode
R10219 N10218 N10219 10
D10219 N10219 0 diode
R10220 N10219 N10220 10
D10220 N10220 0 diode
R10221 N10220 N10221 10
D10221 N10221 0 diode
R10222 N10221 N10222 10
D10222 N10222 0 diode
R10223 N10222 N10223 10
D10223 N10223 0 diode
R10224 N10223 N10224 10
D10224 N10224 0 diode
R10225 N10224 N10225 10
D10225 N10225 0 diode
R10226 N10225 N10226 10
D10226 N10226 0 diode
R10227 N10226 N10227 10
D10227 N10227 0 diode
R10228 N10227 N10228 10
D10228 N10228 0 diode
R10229 N10228 N10229 10
D10229 N10229 0 diode
R10230 N10229 N10230 10
D10230 N10230 0 diode
R10231 N10230 N10231 10
D10231 N10231 0 diode
R10232 N10231 N10232 10
D10232 N10232 0 diode
R10233 N10232 N10233 10
D10233 N10233 0 diode
R10234 N10233 N10234 10
D10234 N10234 0 diode
R10235 N10234 N10235 10
D10235 N10235 0 diode
R10236 N10235 N10236 10
D10236 N10236 0 diode
R10237 N10236 N10237 10
D10237 N10237 0 diode
R10238 N10237 N10238 10
D10238 N10238 0 diode
R10239 N10238 N10239 10
D10239 N10239 0 diode
R10240 N10239 N10240 10
D10240 N10240 0 diode
R10241 N10240 N10241 10
D10241 N10241 0 diode
R10242 N10241 N10242 10
D10242 N10242 0 diode
R10243 N10242 N10243 10
D10243 N10243 0 diode
R10244 N10243 N10244 10
D10244 N10244 0 diode
R10245 N10244 N10245 10
D10245 N10245 0 diode
R10246 N10245 N10246 10
D10246 N10246 0 diode
R10247 N10246 N10247 10
D10247 N10247 0 diode
R10248 N10247 N10248 10
D10248 N10248 0 diode
R10249 N10248 N10249 10
D10249 N10249 0 diode
R10250 N10249 N10250 10
D10250 N10250 0 diode
R10251 N10250 N10251 10
D10251 N10251 0 diode
R10252 N10251 N10252 10
D10252 N10252 0 diode
R10253 N10252 N10253 10
D10253 N10253 0 diode
R10254 N10253 N10254 10
D10254 N10254 0 diode
R10255 N10254 N10255 10
D10255 N10255 0 diode
R10256 N10255 N10256 10
D10256 N10256 0 diode
R10257 N10256 N10257 10
D10257 N10257 0 diode
R10258 N10257 N10258 10
D10258 N10258 0 diode
R10259 N10258 N10259 10
D10259 N10259 0 diode
R10260 N10259 N10260 10
D10260 N10260 0 diode
R10261 N10260 N10261 10
D10261 N10261 0 diode
R10262 N10261 N10262 10
D10262 N10262 0 diode
R10263 N10262 N10263 10
D10263 N10263 0 diode
R10264 N10263 N10264 10
D10264 N10264 0 diode
R10265 N10264 N10265 10
D10265 N10265 0 diode
R10266 N10265 N10266 10
D10266 N10266 0 diode
R10267 N10266 N10267 10
D10267 N10267 0 diode
R10268 N10267 N10268 10
D10268 N10268 0 diode
R10269 N10268 N10269 10
D10269 N10269 0 diode
R10270 N10269 N10270 10
D10270 N10270 0 diode
R10271 N10270 N10271 10
D10271 N10271 0 diode
R10272 N10271 N10272 10
D10272 N10272 0 diode
R10273 N10272 N10273 10
D10273 N10273 0 diode
R10274 N10273 N10274 10
D10274 N10274 0 diode
R10275 N10274 N10275 10
D10275 N10275 0 diode
R10276 N10275 N10276 10
D10276 N10276 0 diode
R10277 N10276 N10277 10
D10277 N10277 0 diode
R10278 N10277 N10278 10
D10278 N10278 0 diode
R10279 N10278 N10279 10
D10279 N10279 0 diode
R10280 N10279 N10280 10
D10280 N10280 0 diode
R10281 N10280 N10281 10
D10281 N10281 0 diode
R10282 N10281 N10282 10
D10282 N10282 0 diode
R10283 N10282 N10283 10
D10283 N10283 0 diode
R10284 N10283 N10284 10
D10284 N10284 0 diode
R10285 N10284 N10285 10
D10285 N10285 0 diode
R10286 N10285 N10286 10
D10286 N10286 0 diode
R10287 N10286 N10287 10
D10287 N10287 0 diode
R10288 N10287 N10288 10
D10288 N10288 0 diode
R10289 N10288 N10289 10
D10289 N10289 0 diode
R10290 N10289 N10290 10
D10290 N10290 0 diode
R10291 N10290 N10291 10
D10291 N10291 0 diode
R10292 N10291 N10292 10
D10292 N10292 0 diode
R10293 N10292 N10293 10
D10293 N10293 0 diode
R10294 N10293 N10294 10
D10294 N10294 0 diode
R10295 N10294 N10295 10
D10295 N10295 0 diode
R10296 N10295 N10296 10
D10296 N10296 0 diode
R10297 N10296 N10297 10
D10297 N10297 0 diode
R10298 N10297 N10298 10
D10298 N10298 0 diode
R10299 N10298 N10299 10
D10299 N10299 0 diode
R10300 N10299 N10300 10
D10300 N10300 0 diode
R10301 N10300 N10301 10
D10301 N10301 0 diode
R10302 N10301 N10302 10
D10302 N10302 0 diode
R10303 N10302 N10303 10
D10303 N10303 0 diode
R10304 N10303 N10304 10
D10304 N10304 0 diode
R10305 N10304 N10305 10
D10305 N10305 0 diode
R10306 N10305 N10306 10
D10306 N10306 0 diode
R10307 N10306 N10307 10
D10307 N10307 0 diode
R10308 N10307 N10308 10
D10308 N10308 0 diode
R10309 N10308 N10309 10
D10309 N10309 0 diode
R10310 N10309 N10310 10
D10310 N10310 0 diode
R10311 N10310 N10311 10
D10311 N10311 0 diode
R10312 N10311 N10312 10
D10312 N10312 0 diode
R10313 N10312 N10313 10
D10313 N10313 0 diode
R10314 N10313 N10314 10
D10314 N10314 0 diode
R10315 N10314 N10315 10
D10315 N10315 0 diode
R10316 N10315 N10316 10
D10316 N10316 0 diode
R10317 N10316 N10317 10
D10317 N10317 0 diode
R10318 N10317 N10318 10
D10318 N10318 0 diode
R10319 N10318 N10319 10
D10319 N10319 0 diode
R10320 N10319 N10320 10
D10320 N10320 0 diode
R10321 N10320 N10321 10
D10321 N10321 0 diode
R10322 N10321 N10322 10
D10322 N10322 0 diode
R10323 N10322 N10323 10
D10323 N10323 0 diode
R10324 N10323 N10324 10
D10324 N10324 0 diode
R10325 N10324 N10325 10
D10325 N10325 0 diode
R10326 N10325 N10326 10
D10326 N10326 0 diode
R10327 N10326 N10327 10
D10327 N10327 0 diode
R10328 N10327 N10328 10
D10328 N10328 0 diode
R10329 N10328 N10329 10
D10329 N10329 0 diode
R10330 N10329 N10330 10
D10330 N10330 0 diode
R10331 N10330 N10331 10
D10331 N10331 0 diode
R10332 N10331 N10332 10
D10332 N10332 0 diode
R10333 N10332 N10333 10
D10333 N10333 0 diode
R10334 N10333 N10334 10
D10334 N10334 0 diode
R10335 N10334 N10335 10
D10335 N10335 0 diode
R10336 N10335 N10336 10
D10336 N10336 0 diode
R10337 N10336 N10337 10
D10337 N10337 0 diode
R10338 N10337 N10338 10
D10338 N10338 0 diode
R10339 N10338 N10339 10
D10339 N10339 0 diode
R10340 N10339 N10340 10
D10340 N10340 0 diode
R10341 N10340 N10341 10
D10341 N10341 0 diode
R10342 N10341 N10342 10
D10342 N10342 0 diode
R10343 N10342 N10343 10
D10343 N10343 0 diode
R10344 N10343 N10344 10
D10344 N10344 0 diode
R10345 N10344 N10345 10
D10345 N10345 0 diode
R10346 N10345 N10346 10
D10346 N10346 0 diode
R10347 N10346 N10347 10
D10347 N10347 0 diode
R10348 N10347 N10348 10
D10348 N10348 0 diode
R10349 N10348 N10349 10
D10349 N10349 0 diode
R10350 N10349 N10350 10
D10350 N10350 0 diode
R10351 N10350 N10351 10
D10351 N10351 0 diode
R10352 N10351 N10352 10
D10352 N10352 0 diode
R10353 N10352 N10353 10
D10353 N10353 0 diode
R10354 N10353 N10354 10
D10354 N10354 0 diode
R10355 N10354 N10355 10
D10355 N10355 0 diode
R10356 N10355 N10356 10
D10356 N10356 0 diode
R10357 N10356 N10357 10
D10357 N10357 0 diode
R10358 N10357 N10358 10
D10358 N10358 0 diode
R10359 N10358 N10359 10
D10359 N10359 0 diode
R10360 N10359 N10360 10
D10360 N10360 0 diode
R10361 N10360 N10361 10
D10361 N10361 0 diode
R10362 N10361 N10362 10
D10362 N10362 0 diode
R10363 N10362 N10363 10
D10363 N10363 0 diode
R10364 N10363 N10364 10
D10364 N10364 0 diode
R10365 N10364 N10365 10
D10365 N10365 0 diode
R10366 N10365 N10366 10
D10366 N10366 0 diode
R10367 N10366 N10367 10
D10367 N10367 0 diode
R10368 N10367 N10368 10
D10368 N10368 0 diode
R10369 N10368 N10369 10
D10369 N10369 0 diode
R10370 N10369 N10370 10
D10370 N10370 0 diode
R10371 N10370 N10371 10
D10371 N10371 0 diode
R10372 N10371 N10372 10
D10372 N10372 0 diode
R10373 N10372 N10373 10
D10373 N10373 0 diode
R10374 N10373 N10374 10
D10374 N10374 0 diode
R10375 N10374 N10375 10
D10375 N10375 0 diode
R10376 N10375 N10376 10
D10376 N10376 0 diode
R10377 N10376 N10377 10
D10377 N10377 0 diode
R10378 N10377 N10378 10
D10378 N10378 0 diode
R10379 N10378 N10379 10
D10379 N10379 0 diode
R10380 N10379 N10380 10
D10380 N10380 0 diode
R10381 N10380 N10381 10
D10381 N10381 0 diode
R10382 N10381 N10382 10
D10382 N10382 0 diode
R10383 N10382 N10383 10
D10383 N10383 0 diode
R10384 N10383 N10384 10
D10384 N10384 0 diode
R10385 N10384 N10385 10
D10385 N10385 0 diode
R10386 N10385 N10386 10
D10386 N10386 0 diode
R10387 N10386 N10387 10
D10387 N10387 0 diode
R10388 N10387 N10388 10
D10388 N10388 0 diode
R10389 N10388 N10389 10
D10389 N10389 0 diode
R10390 N10389 N10390 10
D10390 N10390 0 diode
R10391 N10390 N10391 10
D10391 N10391 0 diode
R10392 N10391 N10392 10
D10392 N10392 0 diode
R10393 N10392 N10393 10
D10393 N10393 0 diode
R10394 N10393 N10394 10
D10394 N10394 0 diode
R10395 N10394 N10395 10
D10395 N10395 0 diode
R10396 N10395 N10396 10
D10396 N10396 0 diode
R10397 N10396 N10397 10
D10397 N10397 0 diode
R10398 N10397 N10398 10
D10398 N10398 0 diode
R10399 N10398 N10399 10
D10399 N10399 0 diode
R10400 N10399 N10400 10
D10400 N10400 0 diode
R10401 N10400 N10401 10
D10401 N10401 0 diode
R10402 N10401 N10402 10
D10402 N10402 0 diode
R10403 N10402 N10403 10
D10403 N10403 0 diode
R10404 N10403 N10404 10
D10404 N10404 0 diode
R10405 N10404 N10405 10
D10405 N10405 0 diode
R10406 N10405 N10406 10
D10406 N10406 0 diode
R10407 N10406 N10407 10
D10407 N10407 0 diode
R10408 N10407 N10408 10
D10408 N10408 0 diode
R10409 N10408 N10409 10
D10409 N10409 0 diode
R10410 N10409 N10410 10
D10410 N10410 0 diode
R10411 N10410 N10411 10
D10411 N10411 0 diode
R10412 N10411 N10412 10
D10412 N10412 0 diode
R10413 N10412 N10413 10
D10413 N10413 0 diode
R10414 N10413 N10414 10
D10414 N10414 0 diode
R10415 N10414 N10415 10
D10415 N10415 0 diode
R10416 N10415 N10416 10
D10416 N10416 0 diode
R10417 N10416 N10417 10
D10417 N10417 0 diode
R10418 N10417 N10418 10
D10418 N10418 0 diode
R10419 N10418 N10419 10
D10419 N10419 0 diode
R10420 N10419 N10420 10
D10420 N10420 0 diode
R10421 N10420 N10421 10
D10421 N10421 0 diode
R10422 N10421 N10422 10
D10422 N10422 0 diode
R10423 N10422 N10423 10
D10423 N10423 0 diode
R10424 N10423 N10424 10
D10424 N10424 0 diode
R10425 N10424 N10425 10
D10425 N10425 0 diode
R10426 N10425 N10426 10
D10426 N10426 0 diode
R10427 N10426 N10427 10
D10427 N10427 0 diode
R10428 N10427 N10428 10
D10428 N10428 0 diode
R10429 N10428 N10429 10
D10429 N10429 0 diode
R10430 N10429 N10430 10
D10430 N10430 0 diode
R10431 N10430 N10431 10
D10431 N10431 0 diode
R10432 N10431 N10432 10
D10432 N10432 0 diode
R10433 N10432 N10433 10
D10433 N10433 0 diode
R10434 N10433 N10434 10
D10434 N10434 0 diode
R10435 N10434 N10435 10
D10435 N10435 0 diode
R10436 N10435 N10436 10
D10436 N10436 0 diode
R10437 N10436 N10437 10
D10437 N10437 0 diode
R10438 N10437 N10438 10
D10438 N10438 0 diode
R10439 N10438 N10439 10
D10439 N10439 0 diode
R10440 N10439 N10440 10
D10440 N10440 0 diode
R10441 N10440 N10441 10
D10441 N10441 0 diode
R10442 N10441 N10442 10
D10442 N10442 0 diode
R10443 N10442 N10443 10
D10443 N10443 0 diode
R10444 N10443 N10444 10
D10444 N10444 0 diode
R10445 N10444 N10445 10
D10445 N10445 0 diode
R10446 N10445 N10446 10
D10446 N10446 0 diode
R10447 N10446 N10447 10
D10447 N10447 0 diode
R10448 N10447 N10448 10
D10448 N10448 0 diode
R10449 N10448 N10449 10
D10449 N10449 0 diode
R10450 N10449 N10450 10
D10450 N10450 0 diode
R10451 N10450 N10451 10
D10451 N10451 0 diode
R10452 N10451 N10452 10
D10452 N10452 0 diode
R10453 N10452 N10453 10
D10453 N10453 0 diode
R10454 N10453 N10454 10
D10454 N10454 0 diode
R10455 N10454 N10455 10
D10455 N10455 0 diode
R10456 N10455 N10456 10
D10456 N10456 0 diode
R10457 N10456 N10457 10
D10457 N10457 0 diode
R10458 N10457 N10458 10
D10458 N10458 0 diode
R10459 N10458 N10459 10
D10459 N10459 0 diode
R10460 N10459 N10460 10
D10460 N10460 0 diode
R10461 N10460 N10461 10
D10461 N10461 0 diode
R10462 N10461 N10462 10
D10462 N10462 0 diode
R10463 N10462 N10463 10
D10463 N10463 0 diode
R10464 N10463 N10464 10
D10464 N10464 0 diode
R10465 N10464 N10465 10
D10465 N10465 0 diode
R10466 N10465 N10466 10
D10466 N10466 0 diode
R10467 N10466 N10467 10
D10467 N10467 0 diode
R10468 N10467 N10468 10
D10468 N10468 0 diode
R10469 N10468 N10469 10
D10469 N10469 0 diode
R10470 N10469 N10470 10
D10470 N10470 0 diode
R10471 N10470 N10471 10
D10471 N10471 0 diode
R10472 N10471 N10472 10
D10472 N10472 0 diode
R10473 N10472 N10473 10
D10473 N10473 0 diode
R10474 N10473 N10474 10
D10474 N10474 0 diode
R10475 N10474 N10475 10
D10475 N10475 0 diode
R10476 N10475 N10476 10
D10476 N10476 0 diode
R10477 N10476 N10477 10
D10477 N10477 0 diode
R10478 N10477 N10478 10
D10478 N10478 0 diode
R10479 N10478 N10479 10
D10479 N10479 0 diode
R10480 N10479 N10480 10
D10480 N10480 0 diode
R10481 N10480 N10481 10
D10481 N10481 0 diode
R10482 N10481 N10482 10
D10482 N10482 0 diode
R10483 N10482 N10483 10
D10483 N10483 0 diode
R10484 N10483 N10484 10
D10484 N10484 0 diode
R10485 N10484 N10485 10
D10485 N10485 0 diode
R10486 N10485 N10486 10
D10486 N10486 0 diode
R10487 N10486 N10487 10
D10487 N10487 0 diode
R10488 N10487 N10488 10
D10488 N10488 0 diode
R10489 N10488 N10489 10
D10489 N10489 0 diode
R10490 N10489 N10490 10
D10490 N10490 0 diode
R10491 N10490 N10491 10
D10491 N10491 0 diode
R10492 N10491 N10492 10
D10492 N10492 0 diode
R10493 N10492 N10493 10
D10493 N10493 0 diode
R10494 N10493 N10494 10
D10494 N10494 0 diode
R10495 N10494 N10495 10
D10495 N10495 0 diode
R10496 N10495 N10496 10
D10496 N10496 0 diode
R10497 N10496 N10497 10
D10497 N10497 0 diode
R10498 N10497 N10498 10
D10498 N10498 0 diode
R10499 N10498 N10499 10
D10499 N10499 0 diode
R10500 N10499 N10500 10
D10500 N10500 0 diode
R10501 N10500 N10501 10
D10501 N10501 0 diode
R10502 N10501 N10502 10
D10502 N10502 0 diode
R10503 N10502 N10503 10
D10503 N10503 0 diode
R10504 N10503 N10504 10
D10504 N10504 0 diode
R10505 N10504 N10505 10
D10505 N10505 0 diode
R10506 N10505 N10506 10
D10506 N10506 0 diode
R10507 N10506 N10507 10
D10507 N10507 0 diode
R10508 N10507 N10508 10
D10508 N10508 0 diode
R10509 N10508 N10509 10
D10509 N10509 0 diode
R10510 N10509 N10510 10
D10510 N10510 0 diode
R10511 N10510 N10511 10
D10511 N10511 0 diode
R10512 N10511 N10512 10
D10512 N10512 0 diode
R10513 N10512 N10513 10
D10513 N10513 0 diode
R10514 N10513 N10514 10
D10514 N10514 0 diode
R10515 N10514 N10515 10
D10515 N10515 0 diode
R10516 N10515 N10516 10
D10516 N10516 0 diode
R10517 N10516 N10517 10
D10517 N10517 0 diode
R10518 N10517 N10518 10
D10518 N10518 0 diode
R10519 N10518 N10519 10
D10519 N10519 0 diode
R10520 N10519 N10520 10
D10520 N10520 0 diode
R10521 N10520 N10521 10
D10521 N10521 0 diode
R10522 N10521 N10522 10
D10522 N10522 0 diode
R10523 N10522 N10523 10
D10523 N10523 0 diode
R10524 N10523 N10524 10
D10524 N10524 0 diode
R10525 N10524 N10525 10
D10525 N10525 0 diode
R10526 N10525 N10526 10
D10526 N10526 0 diode
R10527 N10526 N10527 10
D10527 N10527 0 diode
R10528 N10527 N10528 10
D10528 N10528 0 diode
R10529 N10528 N10529 10
D10529 N10529 0 diode
R10530 N10529 N10530 10
D10530 N10530 0 diode
R10531 N10530 N10531 10
D10531 N10531 0 diode
R10532 N10531 N10532 10
D10532 N10532 0 diode
R10533 N10532 N10533 10
D10533 N10533 0 diode
R10534 N10533 N10534 10
D10534 N10534 0 diode
R10535 N10534 N10535 10
D10535 N10535 0 diode
R10536 N10535 N10536 10
D10536 N10536 0 diode
R10537 N10536 N10537 10
D10537 N10537 0 diode
R10538 N10537 N10538 10
D10538 N10538 0 diode
R10539 N10538 N10539 10
D10539 N10539 0 diode
R10540 N10539 N10540 10
D10540 N10540 0 diode
R10541 N10540 N10541 10
D10541 N10541 0 diode
R10542 N10541 N10542 10
D10542 N10542 0 diode
R10543 N10542 N10543 10
D10543 N10543 0 diode
R10544 N10543 N10544 10
D10544 N10544 0 diode
R10545 N10544 N10545 10
D10545 N10545 0 diode
R10546 N10545 N10546 10
D10546 N10546 0 diode
R10547 N10546 N10547 10
D10547 N10547 0 diode
R10548 N10547 N10548 10
D10548 N10548 0 diode
R10549 N10548 N10549 10
D10549 N10549 0 diode
R10550 N10549 N10550 10
D10550 N10550 0 diode
R10551 N10550 N10551 10
D10551 N10551 0 diode
R10552 N10551 N10552 10
D10552 N10552 0 diode
R10553 N10552 N10553 10
D10553 N10553 0 diode
R10554 N10553 N10554 10
D10554 N10554 0 diode
R10555 N10554 N10555 10
D10555 N10555 0 diode
R10556 N10555 N10556 10
D10556 N10556 0 diode
R10557 N10556 N10557 10
D10557 N10557 0 diode
R10558 N10557 N10558 10
D10558 N10558 0 diode
R10559 N10558 N10559 10
D10559 N10559 0 diode
R10560 N10559 N10560 10
D10560 N10560 0 diode
R10561 N10560 N10561 10
D10561 N10561 0 diode
R10562 N10561 N10562 10
D10562 N10562 0 diode
R10563 N10562 N10563 10
D10563 N10563 0 diode
R10564 N10563 N10564 10
D10564 N10564 0 diode
R10565 N10564 N10565 10
D10565 N10565 0 diode
R10566 N10565 N10566 10
D10566 N10566 0 diode
R10567 N10566 N10567 10
D10567 N10567 0 diode
R10568 N10567 N10568 10
D10568 N10568 0 diode
R10569 N10568 N10569 10
D10569 N10569 0 diode
R10570 N10569 N10570 10
D10570 N10570 0 diode
R10571 N10570 N10571 10
D10571 N10571 0 diode
R10572 N10571 N10572 10
D10572 N10572 0 diode
R10573 N10572 N10573 10
D10573 N10573 0 diode
R10574 N10573 N10574 10
D10574 N10574 0 diode
R10575 N10574 N10575 10
D10575 N10575 0 diode
R10576 N10575 N10576 10
D10576 N10576 0 diode
R10577 N10576 N10577 10
D10577 N10577 0 diode
R10578 N10577 N10578 10
D10578 N10578 0 diode
R10579 N10578 N10579 10
D10579 N10579 0 diode
R10580 N10579 N10580 10
D10580 N10580 0 diode
R10581 N10580 N10581 10
D10581 N10581 0 diode
R10582 N10581 N10582 10
D10582 N10582 0 diode
R10583 N10582 N10583 10
D10583 N10583 0 diode
R10584 N10583 N10584 10
D10584 N10584 0 diode
R10585 N10584 N10585 10
D10585 N10585 0 diode
R10586 N10585 N10586 10
D10586 N10586 0 diode
R10587 N10586 N10587 10
D10587 N10587 0 diode
R10588 N10587 N10588 10
D10588 N10588 0 diode
R10589 N10588 N10589 10
D10589 N10589 0 diode
R10590 N10589 N10590 10
D10590 N10590 0 diode
R10591 N10590 N10591 10
D10591 N10591 0 diode
R10592 N10591 N10592 10
D10592 N10592 0 diode
R10593 N10592 N10593 10
D10593 N10593 0 diode
R10594 N10593 N10594 10
D10594 N10594 0 diode
R10595 N10594 N10595 10
D10595 N10595 0 diode
R10596 N10595 N10596 10
D10596 N10596 0 diode
R10597 N10596 N10597 10
D10597 N10597 0 diode
R10598 N10597 N10598 10
D10598 N10598 0 diode
R10599 N10598 N10599 10
D10599 N10599 0 diode
R10600 N10599 N10600 10
D10600 N10600 0 diode
R10601 N10600 N10601 10
D10601 N10601 0 diode
R10602 N10601 N10602 10
D10602 N10602 0 diode
R10603 N10602 N10603 10
D10603 N10603 0 diode
R10604 N10603 N10604 10
D10604 N10604 0 diode
R10605 N10604 N10605 10
D10605 N10605 0 diode
R10606 N10605 N10606 10
D10606 N10606 0 diode
R10607 N10606 N10607 10
D10607 N10607 0 diode
R10608 N10607 N10608 10
D10608 N10608 0 diode
R10609 N10608 N10609 10
D10609 N10609 0 diode
R10610 N10609 N10610 10
D10610 N10610 0 diode
R10611 N10610 N10611 10
D10611 N10611 0 diode
R10612 N10611 N10612 10
D10612 N10612 0 diode
R10613 N10612 N10613 10
D10613 N10613 0 diode
R10614 N10613 N10614 10
D10614 N10614 0 diode
R10615 N10614 N10615 10
D10615 N10615 0 diode
R10616 N10615 N10616 10
D10616 N10616 0 diode
R10617 N10616 N10617 10
D10617 N10617 0 diode
R10618 N10617 N10618 10
D10618 N10618 0 diode
R10619 N10618 N10619 10
D10619 N10619 0 diode
R10620 N10619 N10620 10
D10620 N10620 0 diode
R10621 N10620 N10621 10
D10621 N10621 0 diode
R10622 N10621 N10622 10
D10622 N10622 0 diode
R10623 N10622 N10623 10
D10623 N10623 0 diode
R10624 N10623 N10624 10
D10624 N10624 0 diode
R10625 N10624 N10625 10
D10625 N10625 0 diode
R10626 N10625 N10626 10
D10626 N10626 0 diode
R10627 N10626 N10627 10
D10627 N10627 0 diode
R10628 N10627 N10628 10
D10628 N10628 0 diode
R10629 N10628 N10629 10
D10629 N10629 0 diode
R10630 N10629 N10630 10
D10630 N10630 0 diode
R10631 N10630 N10631 10
D10631 N10631 0 diode
R10632 N10631 N10632 10
D10632 N10632 0 diode
R10633 N10632 N10633 10
D10633 N10633 0 diode
R10634 N10633 N10634 10
D10634 N10634 0 diode
R10635 N10634 N10635 10
D10635 N10635 0 diode
R10636 N10635 N10636 10
D10636 N10636 0 diode
R10637 N10636 N10637 10
D10637 N10637 0 diode
R10638 N10637 N10638 10
D10638 N10638 0 diode
R10639 N10638 N10639 10
D10639 N10639 0 diode
R10640 N10639 N10640 10
D10640 N10640 0 diode
R10641 N10640 N10641 10
D10641 N10641 0 diode
R10642 N10641 N10642 10
D10642 N10642 0 diode
R10643 N10642 N10643 10
D10643 N10643 0 diode
R10644 N10643 N10644 10
D10644 N10644 0 diode
R10645 N10644 N10645 10
D10645 N10645 0 diode
R10646 N10645 N10646 10
D10646 N10646 0 diode
R10647 N10646 N10647 10
D10647 N10647 0 diode
R10648 N10647 N10648 10
D10648 N10648 0 diode
R10649 N10648 N10649 10
D10649 N10649 0 diode
R10650 N10649 N10650 10
D10650 N10650 0 diode
R10651 N10650 N10651 10
D10651 N10651 0 diode
R10652 N10651 N10652 10
D10652 N10652 0 diode
R10653 N10652 N10653 10
D10653 N10653 0 diode
R10654 N10653 N10654 10
D10654 N10654 0 diode
R10655 N10654 N10655 10
D10655 N10655 0 diode
R10656 N10655 N10656 10
D10656 N10656 0 diode
R10657 N10656 N10657 10
D10657 N10657 0 diode
R10658 N10657 N10658 10
D10658 N10658 0 diode
R10659 N10658 N10659 10
D10659 N10659 0 diode
R10660 N10659 N10660 10
D10660 N10660 0 diode
R10661 N10660 N10661 10
D10661 N10661 0 diode
R10662 N10661 N10662 10
D10662 N10662 0 diode
R10663 N10662 N10663 10
D10663 N10663 0 diode
R10664 N10663 N10664 10
D10664 N10664 0 diode
R10665 N10664 N10665 10
D10665 N10665 0 diode
R10666 N10665 N10666 10
D10666 N10666 0 diode
R10667 N10666 N10667 10
D10667 N10667 0 diode
R10668 N10667 N10668 10
D10668 N10668 0 diode
R10669 N10668 N10669 10
D10669 N10669 0 diode
R10670 N10669 N10670 10
D10670 N10670 0 diode
R10671 N10670 N10671 10
D10671 N10671 0 diode
R10672 N10671 N10672 10
D10672 N10672 0 diode
R10673 N10672 N10673 10
D10673 N10673 0 diode
R10674 N10673 N10674 10
D10674 N10674 0 diode
R10675 N10674 N10675 10
D10675 N10675 0 diode
R10676 N10675 N10676 10
D10676 N10676 0 diode
R10677 N10676 N10677 10
D10677 N10677 0 diode
R10678 N10677 N10678 10
D10678 N10678 0 diode
R10679 N10678 N10679 10
D10679 N10679 0 diode
R10680 N10679 N10680 10
D10680 N10680 0 diode
R10681 N10680 N10681 10
D10681 N10681 0 diode
R10682 N10681 N10682 10
D10682 N10682 0 diode
R10683 N10682 N10683 10
D10683 N10683 0 diode
R10684 N10683 N10684 10
D10684 N10684 0 diode
R10685 N10684 N10685 10
D10685 N10685 0 diode
R10686 N10685 N10686 10
D10686 N10686 0 diode
R10687 N10686 N10687 10
D10687 N10687 0 diode
R10688 N10687 N10688 10
D10688 N10688 0 diode
R10689 N10688 N10689 10
D10689 N10689 0 diode
R10690 N10689 N10690 10
D10690 N10690 0 diode
R10691 N10690 N10691 10
D10691 N10691 0 diode
R10692 N10691 N10692 10
D10692 N10692 0 diode
R10693 N10692 N10693 10
D10693 N10693 0 diode
R10694 N10693 N10694 10
D10694 N10694 0 diode
R10695 N10694 N10695 10
D10695 N10695 0 diode
R10696 N10695 N10696 10
D10696 N10696 0 diode
R10697 N10696 N10697 10
D10697 N10697 0 diode
R10698 N10697 N10698 10
D10698 N10698 0 diode
R10699 N10698 N10699 10
D10699 N10699 0 diode
R10700 N10699 N10700 10
D10700 N10700 0 diode
R10701 N10700 N10701 10
D10701 N10701 0 diode
R10702 N10701 N10702 10
D10702 N10702 0 diode
R10703 N10702 N10703 10
D10703 N10703 0 diode
R10704 N10703 N10704 10
D10704 N10704 0 diode
R10705 N10704 N10705 10
D10705 N10705 0 diode
R10706 N10705 N10706 10
D10706 N10706 0 diode
R10707 N10706 N10707 10
D10707 N10707 0 diode
R10708 N10707 N10708 10
D10708 N10708 0 diode
R10709 N10708 N10709 10
D10709 N10709 0 diode
R10710 N10709 N10710 10
D10710 N10710 0 diode
R10711 N10710 N10711 10
D10711 N10711 0 diode
R10712 N10711 N10712 10
D10712 N10712 0 diode
R10713 N10712 N10713 10
D10713 N10713 0 diode
R10714 N10713 N10714 10
D10714 N10714 0 diode
R10715 N10714 N10715 10
D10715 N10715 0 diode
R10716 N10715 N10716 10
D10716 N10716 0 diode
R10717 N10716 N10717 10
D10717 N10717 0 diode
R10718 N10717 N10718 10
D10718 N10718 0 diode
R10719 N10718 N10719 10
D10719 N10719 0 diode
R10720 N10719 N10720 10
D10720 N10720 0 diode
R10721 N10720 N10721 10
D10721 N10721 0 diode
R10722 N10721 N10722 10
D10722 N10722 0 diode
R10723 N10722 N10723 10
D10723 N10723 0 diode
R10724 N10723 N10724 10
D10724 N10724 0 diode
R10725 N10724 N10725 10
D10725 N10725 0 diode
R10726 N10725 N10726 10
D10726 N10726 0 diode
R10727 N10726 N10727 10
D10727 N10727 0 diode
R10728 N10727 N10728 10
D10728 N10728 0 diode
R10729 N10728 N10729 10
D10729 N10729 0 diode
R10730 N10729 N10730 10
D10730 N10730 0 diode
R10731 N10730 N10731 10
D10731 N10731 0 diode
R10732 N10731 N10732 10
D10732 N10732 0 diode
R10733 N10732 N10733 10
D10733 N10733 0 diode
R10734 N10733 N10734 10
D10734 N10734 0 diode
R10735 N10734 N10735 10
D10735 N10735 0 diode
R10736 N10735 N10736 10
D10736 N10736 0 diode
R10737 N10736 N10737 10
D10737 N10737 0 diode
R10738 N10737 N10738 10
D10738 N10738 0 diode
R10739 N10738 N10739 10
D10739 N10739 0 diode
R10740 N10739 N10740 10
D10740 N10740 0 diode
R10741 N10740 N10741 10
D10741 N10741 0 diode
R10742 N10741 N10742 10
D10742 N10742 0 diode
R10743 N10742 N10743 10
D10743 N10743 0 diode
R10744 N10743 N10744 10
D10744 N10744 0 diode
R10745 N10744 N10745 10
D10745 N10745 0 diode
R10746 N10745 N10746 10
D10746 N10746 0 diode
R10747 N10746 N10747 10
D10747 N10747 0 diode
R10748 N10747 N10748 10
D10748 N10748 0 diode
R10749 N10748 N10749 10
D10749 N10749 0 diode
R10750 N10749 N10750 10
D10750 N10750 0 diode
R10751 N10750 N10751 10
D10751 N10751 0 diode
R10752 N10751 N10752 10
D10752 N10752 0 diode
R10753 N10752 N10753 10
D10753 N10753 0 diode
R10754 N10753 N10754 10
D10754 N10754 0 diode
R10755 N10754 N10755 10
D10755 N10755 0 diode
R10756 N10755 N10756 10
D10756 N10756 0 diode
R10757 N10756 N10757 10
D10757 N10757 0 diode
R10758 N10757 N10758 10
D10758 N10758 0 diode
R10759 N10758 N10759 10
D10759 N10759 0 diode
R10760 N10759 N10760 10
D10760 N10760 0 diode
R10761 N10760 N10761 10
D10761 N10761 0 diode
R10762 N10761 N10762 10
D10762 N10762 0 diode
R10763 N10762 N10763 10
D10763 N10763 0 diode
R10764 N10763 N10764 10
D10764 N10764 0 diode
R10765 N10764 N10765 10
D10765 N10765 0 diode
R10766 N10765 N10766 10
D10766 N10766 0 diode
R10767 N10766 N10767 10
D10767 N10767 0 diode
R10768 N10767 N10768 10
D10768 N10768 0 diode
R10769 N10768 N10769 10
D10769 N10769 0 diode
R10770 N10769 N10770 10
D10770 N10770 0 diode
R10771 N10770 N10771 10
D10771 N10771 0 diode
R10772 N10771 N10772 10
D10772 N10772 0 diode
R10773 N10772 N10773 10
D10773 N10773 0 diode
R10774 N10773 N10774 10
D10774 N10774 0 diode
R10775 N10774 N10775 10
D10775 N10775 0 diode
R10776 N10775 N10776 10
D10776 N10776 0 diode
R10777 N10776 N10777 10
D10777 N10777 0 diode
R10778 N10777 N10778 10
D10778 N10778 0 diode
R10779 N10778 N10779 10
D10779 N10779 0 diode
R10780 N10779 N10780 10
D10780 N10780 0 diode
R10781 N10780 N10781 10
D10781 N10781 0 diode
R10782 N10781 N10782 10
D10782 N10782 0 diode
R10783 N10782 N10783 10
D10783 N10783 0 diode
R10784 N10783 N10784 10
D10784 N10784 0 diode
R10785 N10784 N10785 10
D10785 N10785 0 diode
R10786 N10785 N10786 10
D10786 N10786 0 diode
R10787 N10786 N10787 10
D10787 N10787 0 diode
R10788 N10787 N10788 10
D10788 N10788 0 diode
R10789 N10788 N10789 10
D10789 N10789 0 diode
R10790 N10789 N10790 10
D10790 N10790 0 diode
R10791 N10790 N10791 10
D10791 N10791 0 diode
R10792 N10791 N10792 10
D10792 N10792 0 diode
R10793 N10792 N10793 10
D10793 N10793 0 diode
R10794 N10793 N10794 10
D10794 N10794 0 diode
R10795 N10794 N10795 10
D10795 N10795 0 diode
R10796 N10795 N10796 10
D10796 N10796 0 diode
R10797 N10796 N10797 10
D10797 N10797 0 diode
R10798 N10797 N10798 10
D10798 N10798 0 diode
R10799 N10798 N10799 10
D10799 N10799 0 diode
R10800 N10799 N10800 10
D10800 N10800 0 diode
R10801 N10800 N10801 10
D10801 N10801 0 diode
R10802 N10801 N10802 10
D10802 N10802 0 diode
R10803 N10802 N10803 10
D10803 N10803 0 diode
R10804 N10803 N10804 10
D10804 N10804 0 diode
R10805 N10804 N10805 10
D10805 N10805 0 diode
R10806 N10805 N10806 10
D10806 N10806 0 diode
R10807 N10806 N10807 10
D10807 N10807 0 diode
R10808 N10807 N10808 10
D10808 N10808 0 diode
R10809 N10808 N10809 10
D10809 N10809 0 diode
R10810 N10809 N10810 10
D10810 N10810 0 diode
R10811 N10810 N10811 10
D10811 N10811 0 diode
R10812 N10811 N10812 10
D10812 N10812 0 diode
R10813 N10812 N10813 10
D10813 N10813 0 diode
R10814 N10813 N10814 10
D10814 N10814 0 diode
R10815 N10814 N10815 10
D10815 N10815 0 diode
R10816 N10815 N10816 10
D10816 N10816 0 diode
R10817 N10816 N10817 10
D10817 N10817 0 diode
R10818 N10817 N10818 10
D10818 N10818 0 diode
R10819 N10818 N10819 10
D10819 N10819 0 diode
R10820 N10819 N10820 10
D10820 N10820 0 diode
R10821 N10820 N10821 10
D10821 N10821 0 diode
R10822 N10821 N10822 10
D10822 N10822 0 diode
R10823 N10822 N10823 10
D10823 N10823 0 diode
R10824 N10823 N10824 10
D10824 N10824 0 diode
R10825 N10824 N10825 10
D10825 N10825 0 diode
R10826 N10825 N10826 10
D10826 N10826 0 diode
R10827 N10826 N10827 10
D10827 N10827 0 diode
R10828 N10827 N10828 10
D10828 N10828 0 diode
R10829 N10828 N10829 10
D10829 N10829 0 diode
R10830 N10829 N10830 10
D10830 N10830 0 diode
R10831 N10830 N10831 10
D10831 N10831 0 diode
R10832 N10831 N10832 10
D10832 N10832 0 diode
R10833 N10832 N10833 10
D10833 N10833 0 diode
R10834 N10833 N10834 10
D10834 N10834 0 diode
R10835 N10834 N10835 10
D10835 N10835 0 diode
R10836 N10835 N10836 10
D10836 N10836 0 diode
R10837 N10836 N10837 10
D10837 N10837 0 diode
R10838 N10837 N10838 10
D10838 N10838 0 diode
R10839 N10838 N10839 10
D10839 N10839 0 diode
R10840 N10839 N10840 10
D10840 N10840 0 diode
R10841 N10840 N10841 10
D10841 N10841 0 diode
R10842 N10841 N10842 10
D10842 N10842 0 diode
R10843 N10842 N10843 10
D10843 N10843 0 diode
R10844 N10843 N10844 10
D10844 N10844 0 diode
R10845 N10844 N10845 10
D10845 N10845 0 diode
R10846 N10845 N10846 10
D10846 N10846 0 diode
R10847 N10846 N10847 10
D10847 N10847 0 diode
R10848 N10847 N10848 10
D10848 N10848 0 diode
R10849 N10848 N10849 10
D10849 N10849 0 diode
R10850 N10849 N10850 10
D10850 N10850 0 diode
R10851 N10850 N10851 10
D10851 N10851 0 diode
R10852 N10851 N10852 10
D10852 N10852 0 diode
R10853 N10852 N10853 10
D10853 N10853 0 diode
R10854 N10853 N10854 10
D10854 N10854 0 diode
R10855 N10854 N10855 10
D10855 N10855 0 diode
R10856 N10855 N10856 10
D10856 N10856 0 diode
R10857 N10856 N10857 10
D10857 N10857 0 diode
R10858 N10857 N10858 10
D10858 N10858 0 diode
R10859 N10858 N10859 10
D10859 N10859 0 diode
R10860 N10859 N10860 10
D10860 N10860 0 diode
R10861 N10860 N10861 10
D10861 N10861 0 diode
R10862 N10861 N10862 10
D10862 N10862 0 diode
R10863 N10862 N10863 10
D10863 N10863 0 diode
R10864 N10863 N10864 10
D10864 N10864 0 diode
R10865 N10864 N10865 10
D10865 N10865 0 diode
R10866 N10865 N10866 10
D10866 N10866 0 diode
R10867 N10866 N10867 10
D10867 N10867 0 diode
R10868 N10867 N10868 10
D10868 N10868 0 diode
R10869 N10868 N10869 10
D10869 N10869 0 diode
R10870 N10869 N10870 10
D10870 N10870 0 diode
R10871 N10870 N10871 10
D10871 N10871 0 diode
R10872 N10871 N10872 10
D10872 N10872 0 diode
R10873 N10872 N10873 10
D10873 N10873 0 diode
R10874 N10873 N10874 10
D10874 N10874 0 diode
R10875 N10874 N10875 10
D10875 N10875 0 diode
R10876 N10875 N10876 10
D10876 N10876 0 diode
R10877 N10876 N10877 10
D10877 N10877 0 diode
R10878 N10877 N10878 10
D10878 N10878 0 diode
R10879 N10878 N10879 10
D10879 N10879 0 diode
R10880 N10879 N10880 10
D10880 N10880 0 diode
R10881 N10880 N10881 10
D10881 N10881 0 diode
R10882 N10881 N10882 10
D10882 N10882 0 diode
R10883 N10882 N10883 10
D10883 N10883 0 diode
R10884 N10883 N10884 10
D10884 N10884 0 diode
R10885 N10884 N10885 10
D10885 N10885 0 diode
R10886 N10885 N10886 10
D10886 N10886 0 diode
R10887 N10886 N10887 10
D10887 N10887 0 diode
R10888 N10887 N10888 10
D10888 N10888 0 diode
R10889 N10888 N10889 10
D10889 N10889 0 diode
R10890 N10889 N10890 10
D10890 N10890 0 diode
R10891 N10890 N10891 10
D10891 N10891 0 diode
R10892 N10891 N10892 10
D10892 N10892 0 diode
R10893 N10892 N10893 10
D10893 N10893 0 diode
R10894 N10893 N10894 10
D10894 N10894 0 diode
R10895 N10894 N10895 10
D10895 N10895 0 diode
R10896 N10895 N10896 10
D10896 N10896 0 diode
R10897 N10896 N10897 10
D10897 N10897 0 diode
R10898 N10897 N10898 10
D10898 N10898 0 diode
R10899 N10898 N10899 10
D10899 N10899 0 diode
R10900 N10899 N10900 10
D10900 N10900 0 diode
R10901 N10900 N10901 10
D10901 N10901 0 diode
R10902 N10901 N10902 10
D10902 N10902 0 diode
R10903 N10902 N10903 10
D10903 N10903 0 diode
R10904 N10903 N10904 10
D10904 N10904 0 diode
R10905 N10904 N10905 10
D10905 N10905 0 diode
R10906 N10905 N10906 10
D10906 N10906 0 diode
R10907 N10906 N10907 10
D10907 N10907 0 diode
R10908 N10907 N10908 10
D10908 N10908 0 diode
R10909 N10908 N10909 10
D10909 N10909 0 diode
R10910 N10909 N10910 10
D10910 N10910 0 diode
R10911 N10910 N10911 10
D10911 N10911 0 diode
R10912 N10911 N10912 10
D10912 N10912 0 diode
R10913 N10912 N10913 10
D10913 N10913 0 diode
R10914 N10913 N10914 10
D10914 N10914 0 diode
R10915 N10914 N10915 10
D10915 N10915 0 diode
R10916 N10915 N10916 10
D10916 N10916 0 diode
R10917 N10916 N10917 10
D10917 N10917 0 diode
R10918 N10917 N10918 10
D10918 N10918 0 diode
R10919 N10918 N10919 10
D10919 N10919 0 diode
R10920 N10919 N10920 10
D10920 N10920 0 diode
R10921 N10920 N10921 10
D10921 N10921 0 diode
R10922 N10921 N10922 10
D10922 N10922 0 diode
R10923 N10922 N10923 10
D10923 N10923 0 diode
R10924 N10923 N10924 10
D10924 N10924 0 diode
R10925 N10924 N10925 10
D10925 N10925 0 diode
R10926 N10925 N10926 10
D10926 N10926 0 diode
R10927 N10926 N10927 10
D10927 N10927 0 diode
R10928 N10927 N10928 10
D10928 N10928 0 diode
R10929 N10928 N10929 10
D10929 N10929 0 diode
R10930 N10929 N10930 10
D10930 N10930 0 diode
R10931 N10930 N10931 10
D10931 N10931 0 diode
R10932 N10931 N10932 10
D10932 N10932 0 diode
R10933 N10932 N10933 10
D10933 N10933 0 diode
R10934 N10933 N10934 10
D10934 N10934 0 diode
R10935 N10934 N10935 10
D10935 N10935 0 diode
R10936 N10935 N10936 10
D10936 N10936 0 diode
R10937 N10936 N10937 10
D10937 N10937 0 diode
R10938 N10937 N10938 10
D10938 N10938 0 diode
R10939 N10938 N10939 10
D10939 N10939 0 diode
R10940 N10939 N10940 10
D10940 N10940 0 diode
R10941 N10940 N10941 10
D10941 N10941 0 diode
R10942 N10941 N10942 10
D10942 N10942 0 diode
R10943 N10942 N10943 10
D10943 N10943 0 diode
R10944 N10943 N10944 10
D10944 N10944 0 diode
R10945 N10944 N10945 10
D10945 N10945 0 diode
R10946 N10945 N10946 10
D10946 N10946 0 diode
R10947 N10946 N10947 10
D10947 N10947 0 diode
R10948 N10947 N10948 10
D10948 N10948 0 diode
R10949 N10948 N10949 10
D10949 N10949 0 diode
R10950 N10949 N10950 10
D10950 N10950 0 diode
R10951 N10950 N10951 10
D10951 N10951 0 diode
R10952 N10951 N10952 10
D10952 N10952 0 diode
R10953 N10952 N10953 10
D10953 N10953 0 diode
R10954 N10953 N10954 10
D10954 N10954 0 diode
R10955 N10954 N10955 10
D10955 N10955 0 diode
R10956 N10955 N10956 10
D10956 N10956 0 diode
R10957 N10956 N10957 10
D10957 N10957 0 diode
R10958 N10957 N10958 10
D10958 N10958 0 diode
R10959 N10958 N10959 10
D10959 N10959 0 diode
R10960 N10959 N10960 10
D10960 N10960 0 diode
R10961 N10960 N10961 10
D10961 N10961 0 diode
R10962 N10961 N10962 10
D10962 N10962 0 diode
R10963 N10962 N10963 10
D10963 N10963 0 diode
R10964 N10963 N10964 10
D10964 N10964 0 diode
R10965 N10964 N10965 10
D10965 N10965 0 diode
R10966 N10965 N10966 10
D10966 N10966 0 diode
R10967 N10966 N10967 10
D10967 N10967 0 diode
R10968 N10967 N10968 10
D10968 N10968 0 diode
R10969 N10968 N10969 10
D10969 N10969 0 diode
R10970 N10969 N10970 10
D10970 N10970 0 diode
R10971 N10970 N10971 10
D10971 N10971 0 diode
R10972 N10971 N10972 10
D10972 N10972 0 diode
R10973 N10972 N10973 10
D10973 N10973 0 diode
R10974 N10973 N10974 10
D10974 N10974 0 diode
R10975 N10974 N10975 10
D10975 N10975 0 diode
R10976 N10975 N10976 10
D10976 N10976 0 diode
R10977 N10976 N10977 10
D10977 N10977 0 diode
R10978 N10977 N10978 10
D10978 N10978 0 diode
R10979 N10978 N10979 10
D10979 N10979 0 diode
R10980 N10979 N10980 10
D10980 N10980 0 diode
R10981 N10980 N10981 10
D10981 N10981 0 diode
R10982 N10981 N10982 10
D10982 N10982 0 diode
R10983 N10982 N10983 10
D10983 N10983 0 diode
R10984 N10983 N10984 10
D10984 N10984 0 diode
R10985 N10984 N10985 10
D10985 N10985 0 diode
R10986 N10985 N10986 10
D10986 N10986 0 diode
R10987 N10986 N10987 10
D10987 N10987 0 diode
R10988 N10987 N10988 10
D10988 N10988 0 diode
R10989 N10988 N10989 10
D10989 N10989 0 diode
R10990 N10989 N10990 10
D10990 N10990 0 diode
R10991 N10990 N10991 10
D10991 N10991 0 diode
R10992 N10991 N10992 10
D10992 N10992 0 diode
R10993 N10992 N10993 10
D10993 N10993 0 diode
R10994 N10993 N10994 10
D10994 N10994 0 diode
R10995 N10994 N10995 10
D10995 N10995 0 diode
R10996 N10995 N10996 10
D10996 N10996 0 diode
R10997 N10996 N10997 10
D10997 N10997 0 diode
R10998 N10997 N10998 10
D10998 N10998 0 diode
R10999 N10998 N10999 10
D10999 N10999 0 diode
R11000 N10999 N11000 10
D11000 N11000 0 diode
R11001 N11000 N11001 10
D11001 N11001 0 diode
R11002 N11001 N11002 10
D11002 N11002 0 diode
R11003 N11002 N11003 10
D11003 N11003 0 diode
R11004 N11003 N11004 10
D11004 N11004 0 diode
R11005 N11004 N11005 10
D11005 N11005 0 diode
R11006 N11005 N11006 10
D11006 N11006 0 diode
R11007 N11006 N11007 10
D11007 N11007 0 diode
R11008 N11007 N11008 10
D11008 N11008 0 diode
R11009 N11008 N11009 10
D11009 N11009 0 diode
R11010 N11009 N11010 10
D11010 N11010 0 diode
R11011 N11010 N11011 10
D11011 N11011 0 diode
R11012 N11011 N11012 10
D11012 N11012 0 diode
R11013 N11012 N11013 10
D11013 N11013 0 diode
R11014 N11013 N11014 10
D11014 N11014 0 diode
R11015 N11014 N11015 10
D11015 N11015 0 diode
R11016 N11015 N11016 10
D11016 N11016 0 diode
R11017 N11016 N11017 10
D11017 N11017 0 diode
R11018 N11017 N11018 10
D11018 N11018 0 diode
R11019 N11018 N11019 10
D11019 N11019 0 diode
R11020 N11019 N11020 10
D11020 N11020 0 diode
R11021 N11020 N11021 10
D11021 N11021 0 diode
R11022 N11021 N11022 10
D11022 N11022 0 diode
R11023 N11022 N11023 10
D11023 N11023 0 diode
R11024 N11023 N11024 10
D11024 N11024 0 diode
R11025 N11024 N11025 10
D11025 N11025 0 diode
R11026 N11025 N11026 10
D11026 N11026 0 diode
R11027 N11026 N11027 10
D11027 N11027 0 diode
R11028 N11027 N11028 10
D11028 N11028 0 diode
R11029 N11028 N11029 10
D11029 N11029 0 diode
R11030 N11029 N11030 10
D11030 N11030 0 diode
R11031 N11030 N11031 10
D11031 N11031 0 diode
R11032 N11031 N11032 10
D11032 N11032 0 diode
R11033 N11032 N11033 10
D11033 N11033 0 diode
R11034 N11033 N11034 10
D11034 N11034 0 diode
R11035 N11034 N11035 10
D11035 N11035 0 diode
R11036 N11035 N11036 10
D11036 N11036 0 diode
R11037 N11036 N11037 10
D11037 N11037 0 diode
R11038 N11037 N11038 10
D11038 N11038 0 diode
R11039 N11038 N11039 10
D11039 N11039 0 diode
R11040 N11039 N11040 10
D11040 N11040 0 diode
R11041 N11040 N11041 10
D11041 N11041 0 diode
R11042 N11041 N11042 10
D11042 N11042 0 diode
R11043 N11042 N11043 10
D11043 N11043 0 diode
R11044 N11043 N11044 10
D11044 N11044 0 diode
R11045 N11044 N11045 10
D11045 N11045 0 diode
R11046 N11045 N11046 10
D11046 N11046 0 diode
R11047 N11046 N11047 10
D11047 N11047 0 diode
R11048 N11047 N11048 10
D11048 N11048 0 diode
R11049 N11048 N11049 10
D11049 N11049 0 diode
R11050 N11049 N11050 10
D11050 N11050 0 diode
R11051 N11050 N11051 10
D11051 N11051 0 diode
R11052 N11051 N11052 10
D11052 N11052 0 diode
R11053 N11052 N11053 10
D11053 N11053 0 diode
R11054 N11053 N11054 10
D11054 N11054 0 diode
R11055 N11054 N11055 10
D11055 N11055 0 diode
R11056 N11055 N11056 10
D11056 N11056 0 diode
R11057 N11056 N11057 10
D11057 N11057 0 diode
R11058 N11057 N11058 10
D11058 N11058 0 diode
R11059 N11058 N11059 10
D11059 N11059 0 diode
R11060 N11059 N11060 10
D11060 N11060 0 diode
R11061 N11060 N11061 10
D11061 N11061 0 diode
R11062 N11061 N11062 10
D11062 N11062 0 diode
R11063 N11062 N11063 10
D11063 N11063 0 diode
R11064 N11063 N11064 10
D11064 N11064 0 diode
R11065 N11064 N11065 10
D11065 N11065 0 diode
R11066 N11065 N11066 10
D11066 N11066 0 diode
R11067 N11066 N11067 10
D11067 N11067 0 diode
R11068 N11067 N11068 10
D11068 N11068 0 diode
R11069 N11068 N11069 10
D11069 N11069 0 diode
R11070 N11069 N11070 10
D11070 N11070 0 diode
R11071 N11070 N11071 10
D11071 N11071 0 diode
R11072 N11071 N11072 10
D11072 N11072 0 diode
R11073 N11072 N11073 10
D11073 N11073 0 diode
R11074 N11073 N11074 10
D11074 N11074 0 diode
R11075 N11074 N11075 10
D11075 N11075 0 diode
R11076 N11075 N11076 10
D11076 N11076 0 diode
R11077 N11076 N11077 10
D11077 N11077 0 diode
R11078 N11077 N11078 10
D11078 N11078 0 diode
R11079 N11078 N11079 10
D11079 N11079 0 diode
R11080 N11079 N11080 10
D11080 N11080 0 diode
R11081 N11080 N11081 10
D11081 N11081 0 diode
R11082 N11081 N11082 10
D11082 N11082 0 diode
R11083 N11082 N11083 10
D11083 N11083 0 diode
R11084 N11083 N11084 10
D11084 N11084 0 diode
R11085 N11084 N11085 10
D11085 N11085 0 diode
R11086 N11085 N11086 10
D11086 N11086 0 diode
R11087 N11086 N11087 10
D11087 N11087 0 diode
R11088 N11087 N11088 10
D11088 N11088 0 diode
R11089 N11088 N11089 10
D11089 N11089 0 diode
R11090 N11089 N11090 10
D11090 N11090 0 diode
R11091 N11090 N11091 10
D11091 N11091 0 diode
R11092 N11091 N11092 10
D11092 N11092 0 diode
R11093 N11092 N11093 10
D11093 N11093 0 diode
R11094 N11093 N11094 10
D11094 N11094 0 diode
R11095 N11094 N11095 10
D11095 N11095 0 diode
R11096 N11095 N11096 10
D11096 N11096 0 diode
R11097 N11096 N11097 10
D11097 N11097 0 diode
R11098 N11097 N11098 10
D11098 N11098 0 diode
R11099 N11098 N11099 10
D11099 N11099 0 diode
R11100 N11099 N11100 10
D11100 N11100 0 diode
R11101 N11100 N11101 10
D11101 N11101 0 diode
R11102 N11101 N11102 10
D11102 N11102 0 diode
R11103 N11102 N11103 10
D11103 N11103 0 diode
R11104 N11103 N11104 10
D11104 N11104 0 diode
R11105 N11104 N11105 10
D11105 N11105 0 diode
R11106 N11105 N11106 10
D11106 N11106 0 diode
R11107 N11106 N11107 10
D11107 N11107 0 diode
R11108 N11107 N11108 10
D11108 N11108 0 diode
R11109 N11108 N11109 10
D11109 N11109 0 diode
R11110 N11109 N11110 10
D11110 N11110 0 diode
R11111 N11110 N11111 10
D11111 N11111 0 diode
R11112 N11111 N11112 10
D11112 N11112 0 diode
R11113 N11112 N11113 10
D11113 N11113 0 diode
R11114 N11113 N11114 10
D11114 N11114 0 diode
R11115 N11114 N11115 10
D11115 N11115 0 diode
R11116 N11115 N11116 10
D11116 N11116 0 diode
R11117 N11116 N11117 10
D11117 N11117 0 diode
R11118 N11117 N11118 10
D11118 N11118 0 diode
R11119 N11118 N11119 10
D11119 N11119 0 diode
R11120 N11119 N11120 10
D11120 N11120 0 diode
R11121 N11120 N11121 10
D11121 N11121 0 diode
R11122 N11121 N11122 10
D11122 N11122 0 diode
R11123 N11122 N11123 10
D11123 N11123 0 diode
R11124 N11123 N11124 10
D11124 N11124 0 diode
R11125 N11124 N11125 10
D11125 N11125 0 diode
R11126 N11125 N11126 10
D11126 N11126 0 diode
R11127 N11126 N11127 10
D11127 N11127 0 diode
R11128 N11127 N11128 10
D11128 N11128 0 diode
R11129 N11128 N11129 10
D11129 N11129 0 diode
R11130 N11129 N11130 10
D11130 N11130 0 diode
R11131 N11130 N11131 10
D11131 N11131 0 diode
R11132 N11131 N11132 10
D11132 N11132 0 diode
R11133 N11132 N11133 10
D11133 N11133 0 diode
R11134 N11133 N11134 10
D11134 N11134 0 diode
R11135 N11134 N11135 10
D11135 N11135 0 diode
R11136 N11135 N11136 10
D11136 N11136 0 diode
R11137 N11136 N11137 10
D11137 N11137 0 diode
R11138 N11137 N11138 10
D11138 N11138 0 diode
R11139 N11138 N11139 10
D11139 N11139 0 diode
R11140 N11139 N11140 10
D11140 N11140 0 diode
R11141 N11140 N11141 10
D11141 N11141 0 diode
R11142 N11141 N11142 10
D11142 N11142 0 diode
R11143 N11142 N11143 10
D11143 N11143 0 diode
R11144 N11143 N11144 10
D11144 N11144 0 diode
R11145 N11144 N11145 10
D11145 N11145 0 diode
R11146 N11145 N11146 10
D11146 N11146 0 diode
R11147 N11146 N11147 10
D11147 N11147 0 diode
R11148 N11147 N11148 10
D11148 N11148 0 diode
R11149 N11148 N11149 10
D11149 N11149 0 diode
R11150 N11149 N11150 10
D11150 N11150 0 diode
R11151 N11150 N11151 10
D11151 N11151 0 diode
R11152 N11151 N11152 10
D11152 N11152 0 diode
R11153 N11152 N11153 10
D11153 N11153 0 diode
R11154 N11153 N11154 10
D11154 N11154 0 diode
R11155 N11154 N11155 10
D11155 N11155 0 diode
R11156 N11155 N11156 10
D11156 N11156 0 diode
R11157 N11156 N11157 10
D11157 N11157 0 diode
R11158 N11157 N11158 10
D11158 N11158 0 diode
R11159 N11158 N11159 10
D11159 N11159 0 diode
R11160 N11159 N11160 10
D11160 N11160 0 diode
R11161 N11160 N11161 10
D11161 N11161 0 diode
R11162 N11161 N11162 10
D11162 N11162 0 diode
R11163 N11162 N11163 10
D11163 N11163 0 diode
R11164 N11163 N11164 10
D11164 N11164 0 diode
R11165 N11164 N11165 10
D11165 N11165 0 diode
R11166 N11165 N11166 10
D11166 N11166 0 diode
R11167 N11166 N11167 10
D11167 N11167 0 diode
R11168 N11167 N11168 10
D11168 N11168 0 diode
R11169 N11168 N11169 10
D11169 N11169 0 diode
R11170 N11169 N11170 10
D11170 N11170 0 diode
R11171 N11170 N11171 10
D11171 N11171 0 diode
R11172 N11171 N11172 10
D11172 N11172 0 diode
R11173 N11172 N11173 10
D11173 N11173 0 diode
R11174 N11173 N11174 10
D11174 N11174 0 diode
R11175 N11174 N11175 10
D11175 N11175 0 diode
R11176 N11175 N11176 10
D11176 N11176 0 diode
R11177 N11176 N11177 10
D11177 N11177 0 diode
R11178 N11177 N11178 10
D11178 N11178 0 diode
R11179 N11178 N11179 10
D11179 N11179 0 diode
R11180 N11179 N11180 10
D11180 N11180 0 diode
R11181 N11180 N11181 10
D11181 N11181 0 diode
R11182 N11181 N11182 10
D11182 N11182 0 diode
R11183 N11182 N11183 10
D11183 N11183 0 diode
R11184 N11183 N11184 10
D11184 N11184 0 diode
R11185 N11184 N11185 10
D11185 N11185 0 diode
R11186 N11185 N11186 10
D11186 N11186 0 diode
R11187 N11186 N11187 10
D11187 N11187 0 diode
R11188 N11187 N11188 10
D11188 N11188 0 diode
R11189 N11188 N11189 10
D11189 N11189 0 diode
R11190 N11189 N11190 10
D11190 N11190 0 diode
R11191 N11190 N11191 10
D11191 N11191 0 diode
R11192 N11191 N11192 10
D11192 N11192 0 diode
R11193 N11192 N11193 10
D11193 N11193 0 diode
R11194 N11193 N11194 10
D11194 N11194 0 diode
R11195 N11194 N11195 10
D11195 N11195 0 diode
R11196 N11195 N11196 10
D11196 N11196 0 diode
R11197 N11196 N11197 10
D11197 N11197 0 diode
R11198 N11197 N11198 10
D11198 N11198 0 diode
R11199 N11198 N11199 10
D11199 N11199 0 diode
R11200 N11199 N11200 10
D11200 N11200 0 diode
R11201 N11200 N11201 10
D11201 N11201 0 diode
R11202 N11201 N11202 10
D11202 N11202 0 diode
R11203 N11202 N11203 10
D11203 N11203 0 diode
R11204 N11203 N11204 10
D11204 N11204 0 diode
R11205 N11204 N11205 10
D11205 N11205 0 diode
R11206 N11205 N11206 10
D11206 N11206 0 diode
R11207 N11206 N11207 10
D11207 N11207 0 diode
R11208 N11207 N11208 10
D11208 N11208 0 diode
R11209 N11208 N11209 10
D11209 N11209 0 diode
R11210 N11209 N11210 10
D11210 N11210 0 diode
R11211 N11210 N11211 10
D11211 N11211 0 diode
R11212 N11211 N11212 10
D11212 N11212 0 diode
R11213 N11212 N11213 10
D11213 N11213 0 diode
R11214 N11213 N11214 10
D11214 N11214 0 diode
R11215 N11214 N11215 10
D11215 N11215 0 diode
R11216 N11215 N11216 10
D11216 N11216 0 diode
R11217 N11216 N11217 10
D11217 N11217 0 diode
R11218 N11217 N11218 10
D11218 N11218 0 diode
R11219 N11218 N11219 10
D11219 N11219 0 diode
R11220 N11219 N11220 10
D11220 N11220 0 diode
R11221 N11220 N11221 10
D11221 N11221 0 diode
R11222 N11221 N11222 10
D11222 N11222 0 diode
R11223 N11222 N11223 10
D11223 N11223 0 diode
R11224 N11223 N11224 10
D11224 N11224 0 diode
R11225 N11224 N11225 10
D11225 N11225 0 diode
R11226 N11225 N11226 10
D11226 N11226 0 diode
R11227 N11226 N11227 10
D11227 N11227 0 diode
R11228 N11227 N11228 10
D11228 N11228 0 diode
R11229 N11228 N11229 10
D11229 N11229 0 diode
R11230 N11229 N11230 10
D11230 N11230 0 diode
R11231 N11230 N11231 10
D11231 N11231 0 diode
R11232 N11231 N11232 10
D11232 N11232 0 diode
R11233 N11232 N11233 10
D11233 N11233 0 diode
R11234 N11233 N11234 10
D11234 N11234 0 diode
R11235 N11234 N11235 10
D11235 N11235 0 diode
R11236 N11235 N11236 10
D11236 N11236 0 diode
R11237 N11236 N11237 10
D11237 N11237 0 diode
R11238 N11237 N11238 10
D11238 N11238 0 diode
R11239 N11238 N11239 10
D11239 N11239 0 diode
R11240 N11239 N11240 10
D11240 N11240 0 diode
R11241 N11240 N11241 10
D11241 N11241 0 diode
R11242 N11241 N11242 10
D11242 N11242 0 diode
R11243 N11242 N11243 10
D11243 N11243 0 diode
R11244 N11243 N11244 10
D11244 N11244 0 diode
R11245 N11244 N11245 10
D11245 N11245 0 diode
R11246 N11245 N11246 10
D11246 N11246 0 diode
R11247 N11246 N11247 10
D11247 N11247 0 diode
R11248 N11247 N11248 10
D11248 N11248 0 diode
R11249 N11248 N11249 10
D11249 N11249 0 diode
R11250 N11249 N11250 10
D11250 N11250 0 diode
R11251 N11250 N11251 10
D11251 N11251 0 diode
R11252 N11251 N11252 10
D11252 N11252 0 diode
R11253 N11252 N11253 10
D11253 N11253 0 diode
R11254 N11253 N11254 10
D11254 N11254 0 diode
R11255 N11254 N11255 10
D11255 N11255 0 diode
R11256 N11255 N11256 10
D11256 N11256 0 diode
R11257 N11256 N11257 10
D11257 N11257 0 diode
R11258 N11257 N11258 10
D11258 N11258 0 diode
R11259 N11258 N11259 10
D11259 N11259 0 diode
R11260 N11259 N11260 10
D11260 N11260 0 diode
R11261 N11260 N11261 10
D11261 N11261 0 diode
R11262 N11261 N11262 10
D11262 N11262 0 diode
R11263 N11262 N11263 10
D11263 N11263 0 diode
R11264 N11263 N11264 10
D11264 N11264 0 diode
R11265 N11264 N11265 10
D11265 N11265 0 diode
R11266 N11265 N11266 10
D11266 N11266 0 diode
R11267 N11266 N11267 10
D11267 N11267 0 diode
R11268 N11267 N11268 10
D11268 N11268 0 diode
R11269 N11268 N11269 10
D11269 N11269 0 diode
R11270 N11269 N11270 10
D11270 N11270 0 diode
R11271 N11270 N11271 10
D11271 N11271 0 diode
R11272 N11271 N11272 10
D11272 N11272 0 diode
R11273 N11272 N11273 10
D11273 N11273 0 diode
R11274 N11273 N11274 10
D11274 N11274 0 diode
R11275 N11274 N11275 10
D11275 N11275 0 diode
R11276 N11275 N11276 10
D11276 N11276 0 diode
R11277 N11276 N11277 10
D11277 N11277 0 diode
R11278 N11277 N11278 10
D11278 N11278 0 diode
R11279 N11278 N11279 10
D11279 N11279 0 diode
R11280 N11279 N11280 10
D11280 N11280 0 diode
R11281 N11280 N11281 10
D11281 N11281 0 diode
R11282 N11281 N11282 10
D11282 N11282 0 diode
R11283 N11282 N11283 10
D11283 N11283 0 diode
R11284 N11283 N11284 10
D11284 N11284 0 diode
R11285 N11284 N11285 10
D11285 N11285 0 diode
R11286 N11285 N11286 10
D11286 N11286 0 diode
R11287 N11286 N11287 10
D11287 N11287 0 diode
R11288 N11287 N11288 10
D11288 N11288 0 diode
R11289 N11288 N11289 10
D11289 N11289 0 diode
R11290 N11289 N11290 10
D11290 N11290 0 diode
R11291 N11290 N11291 10
D11291 N11291 0 diode
R11292 N11291 N11292 10
D11292 N11292 0 diode
R11293 N11292 N11293 10
D11293 N11293 0 diode
R11294 N11293 N11294 10
D11294 N11294 0 diode
R11295 N11294 N11295 10
D11295 N11295 0 diode
R11296 N11295 N11296 10
D11296 N11296 0 diode
R11297 N11296 N11297 10
D11297 N11297 0 diode
R11298 N11297 N11298 10
D11298 N11298 0 diode
R11299 N11298 N11299 10
D11299 N11299 0 diode
R11300 N11299 N11300 10
D11300 N11300 0 diode
R11301 N11300 N11301 10
D11301 N11301 0 diode
R11302 N11301 N11302 10
D11302 N11302 0 diode
R11303 N11302 N11303 10
D11303 N11303 0 diode
R11304 N11303 N11304 10
D11304 N11304 0 diode
R11305 N11304 N11305 10
D11305 N11305 0 diode
R11306 N11305 N11306 10
D11306 N11306 0 diode
R11307 N11306 N11307 10
D11307 N11307 0 diode
R11308 N11307 N11308 10
D11308 N11308 0 diode
R11309 N11308 N11309 10
D11309 N11309 0 diode
R11310 N11309 N11310 10
D11310 N11310 0 diode
R11311 N11310 N11311 10
D11311 N11311 0 diode
R11312 N11311 N11312 10
D11312 N11312 0 diode
R11313 N11312 N11313 10
D11313 N11313 0 diode
R11314 N11313 N11314 10
D11314 N11314 0 diode
R11315 N11314 N11315 10
D11315 N11315 0 diode
R11316 N11315 N11316 10
D11316 N11316 0 diode
R11317 N11316 N11317 10
D11317 N11317 0 diode
R11318 N11317 N11318 10
D11318 N11318 0 diode
R11319 N11318 N11319 10
D11319 N11319 0 diode
R11320 N11319 N11320 10
D11320 N11320 0 diode
R11321 N11320 N11321 10
D11321 N11321 0 diode
R11322 N11321 N11322 10
D11322 N11322 0 diode
R11323 N11322 N11323 10
D11323 N11323 0 diode
R11324 N11323 N11324 10
D11324 N11324 0 diode
R11325 N11324 N11325 10
D11325 N11325 0 diode
R11326 N11325 N11326 10
D11326 N11326 0 diode
R11327 N11326 N11327 10
D11327 N11327 0 diode
R11328 N11327 N11328 10
D11328 N11328 0 diode
R11329 N11328 N11329 10
D11329 N11329 0 diode
R11330 N11329 N11330 10
D11330 N11330 0 diode
R11331 N11330 N11331 10
D11331 N11331 0 diode
R11332 N11331 N11332 10
D11332 N11332 0 diode
R11333 N11332 N11333 10
D11333 N11333 0 diode
R11334 N11333 N11334 10
D11334 N11334 0 diode
R11335 N11334 N11335 10
D11335 N11335 0 diode
R11336 N11335 N11336 10
D11336 N11336 0 diode
R11337 N11336 N11337 10
D11337 N11337 0 diode
R11338 N11337 N11338 10
D11338 N11338 0 diode
R11339 N11338 N11339 10
D11339 N11339 0 diode
R11340 N11339 N11340 10
D11340 N11340 0 diode
R11341 N11340 N11341 10
D11341 N11341 0 diode
R11342 N11341 N11342 10
D11342 N11342 0 diode
R11343 N11342 N11343 10
D11343 N11343 0 diode
R11344 N11343 N11344 10
D11344 N11344 0 diode
R11345 N11344 N11345 10
D11345 N11345 0 diode
R11346 N11345 N11346 10
D11346 N11346 0 diode
R11347 N11346 N11347 10
D11347 N11347 0 diode
R11348 N11347 N11348 10
D11348 N11348 0 diode
R11349 N11348 N11349 10
D11349 N11349 0 diode
R11350 N11349 N11350 10
D11350 N11350 0 diode
R11351 N11350 N11351 10
D11351 N11351 0 diode
R11352 N11351 N11352 10
D11352 N11352 0 diode
R11353 N11352 N11353 10
D11353 N11353 0 diode
R11354 N11353 N11354 10
D11354 N11354 0 diode
R11355 N11354 N11355 10
D11355 N11355 0 diode
R11356 N11355 N11356 10
D11356 N11356 0 diode
R11357 N11356 N11357 10
D11357 N11357 0 diode
R11358 N11357 N11358 10
D11358 N11358 0 diode
R11359 N11358 N11359 10
D11359 N11359 0 diode
R11360 N11359 N11360 10
D11360 N11360 0 diode
R11361 N11360 N11361 10
D11361 N11361 0 diode
R11362 N11361 N11362 10
D11362 N11362 0 diode
R11363 N11362 N11363 10
D11363 N11363 0 diode
R11364 N11363 N11364 10
D11364 N11364 0 diode
R11365 N11364 N11365 10
D11365 N11365 0 diode
R11366 N11365 N11366 10
D11366 N11366 0 diode
R11367 N11366 N11367 10
D11367 N11367 0 diode
R11368 N11367 N11368 10
D11368 N11368 0 diode
R11369 N11368 N11369 10
D11369 N11369 0 diode
R11370 N11369 N11370 10
D11370 N11370 0 diode
R11371 N11370 N11371 10
D11371 N11371 0 diode
R11372 N11371 N11372 10
D11372 N11372 0 diode
R11373 N11372 N11373 10
D11373 N11373 0 diode
R11374 N11373 N11374 10
D11374 N11374 0 diode
R11375 N11374 N11375 10
D11375 N11375 0 diode
R11376 N11375 N11376 10
D11376 N11376 0 diode
R11377 N11376 N11377 10
D11377 N11377 0 diode
R11378 N11377 N11378 10
D11378 N11378 0 diode
R11379 N11378 N11379 10
D11379 N11379 0 diode
R11380 N11379 N11380 10
D11380 N11380 0 diode
R11381 N11380 N11381 10
D11381 N11381 0 diode
R11382 N11381 N11382 10
D11382 N11382 0 diode
R11383 N11382 N11383 10
D11383 N11383 0 diode
R11384 N11383 N11384 10
D11384 N11384 0 diode
R11385 N11384 N11385 10
D11385 N11385 0 diode
R11386 N11385 N11386 10
D11386 N11386 0 diode
R11387 N11386 N11387 10
D11387 N11387 0 diode
R11388 N11387 N11388 10
D11388 N11388 0 diode
R11389 N11388 N11389 10
D11389 N11389 0 diode
R11390 N11389 N11390 10
D11390 N11390 0 diode
R11391 N11390 N11391 10
D11391 N11391 0 diode
R11392 N11391 N11392 10
D11392 N11392 0 diode
R11393 N11392 N11393 10
D11393 N11393 0 diode
R11394 N11393 N11394 10
D11394 N11394 0 diode
R11395 N11394 N11395 10
D11395 N11395 0 diode
R11396 N11395 N11396 10
D11396 N11396 0 diode
R11397 N11396 N11397 10
D11397 N11397 0 diode
R11398 N11397 N11398 10
D11398 N11398 0 diode
R11399 N11398 N11399 10
D11399 N11399 0 diode
R11400 N11399 N11400 10
D11400 N11400 0 diode
R11401 N11400 N11401 10
D11401 N11401 0 diode
R11402 N11401 N11402 10
D11402 N11402 0 diode
R11403 N11402 N11403 10
D11403 N11403 0 diode
R11404 N11403 N11404 10
D11404 N11404 0 diode
R11405 N11404 N11405 10
D11405 N11405 0 diode
R11406 N11405 N11406 10
D11406 N11406 0 diode
R11407 N11406 N11407 10
D11407 N11407 0 diode
R11408 N11407 N11408 10
D11408 N11408 0 diode
R11409 N11408 N11409 10
D11409 N11409 0 diode
R11410 N11409 N11410 10
D11410 N11410 0 diode
R11411 N11410 N11411 10
D11411 N11411 0 diode
R11412 N11411 N11412 10
D11412 N11412 0 diode
R11413 N11412 N11413 10
D11413 N11413 0 diode
R11414 N11413 N11414 10
D11414 N11414 0 diode
R11415 N11414 N11415 10
D11415 N11415 0 diode
R11416 N11415 N11416 10
D11416 N11416 0 diode
R11417 N11416 N11417 10
D11417 N11417 0 diode
R11418 N11417 N11418 10
D11418 N11418 0 diode
R11419 N11418 N11419 10
D11419 N11419 0 diode
R11420 N11419 N11420 10
D11420 N11420 0 diode
R11421 N11420 N11421 10
D11421 N11421 0 diode
R11422 N11421 N11422 10
D11422 N11422 0 diode
R11423 N11422 N11423 10
D11423 N11423 0 diode
R11424 N11423 N11424 10
D11424 N11424 0 diode
R11425 N11424 N11425 10
D11425 N11425 0 diode
R11426 N11425 N11426 10
D11426 N11426 0 diode
R11427 N11426 N11427 10
D11427 N11427 0 diode
R11428 N11427 N11428 10
D11428 N11428 0 diode
R11429 N11428 N11429 10
D11429 N11429 0 diode
R11430 N11429 N11430 10
D11430 N11430 0 diode
R11431 N11430 N11431 10
D11431 N11431 0 diode
R11432 N11431 N11432 10
D11432 N11432 0 diode
R11433 N11432 N11433 10
D11433 N11433 0 diode
R11434 N11433 N11434 10
D11434 N11434 0 diode
R11435 N11434 N11435 10
D11435 N11435 0 diode
R11436 N11435 N11436 10
D11436 N11436 0 diode
R11437 N11436 N11437 10
D11437 N11437 0 diode
R11438 N11437 N11438 10
D11438 N11438 0 diode
R11439 N11438 N11439 10
D11439 N11439 0 diode
R11440 N11439 N11440 10
D11440 N11440 0 diode
R11441 N11440 N11441 10
D11441 N11441 0 diode
R11442 N11441 N11442 10
D11442 N11442 0 diode
R11443 N11442 N11443 10
D11443 N11443 0 diode
R11444 N11443 N11444 10
D11444 N11444 0 diode
R11445 N11444 N11445 10
D11445 N11445 0 diode
R11446 N11445 N11446 10
D11446 N11446 0 diode
R11447 N11446 N11447 10
D11447 N11447 0 diode
R11448 N11447 N11448 10
D11448 N11448 0 diode
R11449 N11448 N11449 10
D11449 N11449 0 diode
R11450 N11449 N11450 10
D11450 N11450 0 diode
R11451 N11450 N11451 10
D11451 N11451 0 diode
R11452 N11451 N11452 10
D11452 N11452 0 diode
R11453 N11452 N11453 10
D11453 N11453 0 diode
R11454 N11453 N11454 10
D11454 N11454 0 diode
R11455 N11454 N11455 10
D11455 N11455 0 diode
R11456 N11455 N11456 10
D11456 N11456 0 diode
R11457 N11456 N11457 10
D11457 N11457 0 diode
R11458 N11457 N11458 10
D11458 N11458 0 diode
R11459 N11458 N11459 10
D11459 N11459 0 diode
R11460 N11459 N11460 10
D11460 N11460 0 diode
R11461 N11460 N11461 10
D11461 N11461 0 diode
R11462 N11461 N11462 10
D11462 N11462 0 diode
R11463 N11462 N11463 10
D11463 N11463 0 diode
R11464 N11463 N11464 10
D11464 N11464 0 diode
R11465 N11464 N11465 10
D11465 N11465 0 diode
R11466 N11465 N11466 10
D11466 N11466 0 diode
R11467 N11466 N11467 10
D11467 N11467 0 diode
R11468 N11467 N11468 10
D11468 N11468 0 diode
R11469 N11468 N11469 10
D11469 N11469 0 diode
R11470 N11469 N11470 10
D11470 N11470 0 diode
R11471 N11470 N11471 10
D11471 N11471 0 diode
R11472 N11471 N11472 10
D11472 N11472 0 diode
R11473 N11472 N11473 10
D11473 N11473 0 diode
R11474 N11473 N11474 10
D11474 N11474 0 diode
R11475 N11474 N11475 10
D11475 N11475 0 diode
R11476 N11475 N11476 10
D11476 N11476 0 diode
R11477 N11476 N11477 10
D11477 N11477 0 diode
R11478 N11477 N11478 10
D11478 N11478 0 diode
R11479 N11478 N11479 10
D11479 N11479 0 diode
R11480 N11479 N11480 10
D11480 N11480 0 diode
R11481 N11480 N11481 10
D11481 N11481 0 diode
R11482 N11481 N11482 10
D11482 N11482 0 diode
R11483 N11482 N11483 10
D11483 N11483 0 diode
R11484 N11483 N11484 10
D11484 N11484 0 diode
R11485 N11484 N11485 10
D11485 N11485 0 diode
R11486 N11485 N11486 10
D11486 N11486 0 diode
R11487 N11486 N11487 10
D11487 N11487 0 diode
R11488 N11487 N11488 10
D11488 N11488 0 diode
R11489 N11488 N11489 10
D11489 N11489 0 diode
R11490 N11489 N11490 10
D11490 N11490 0 diode
R11491 N11490 N11491 10
D11491 N11491 0 diode
R11492 N11491 N11492 10
D11492 N11492 0 diode
R11493 N11492 N11493 10
D11493 N11493 0 diode
R11494 N11493 N11494 10
D11494 N11494 0 diode
R11495 N11494 N11495 10
D11495 N11495 0 diode
R11496 N11495 N11496 10
D11496 N11496 0 diode
R11497 N11496 N11497 10
D11497 N11497 0 diode
R11498 N11497 N11498 10
D11498 N11498 0 diode
R11499 N11498 N11499 10
D11499 N11499 0 diode
R11500 N11499 N11500 10
D11500 N11500 0 diode
R11501 N11500 N11501 10
D11501 N11501 0 diode
R11502 N11501 N11502 10
D11502 N11502 0 diode
R11503 N11502 N11503 10
D11503 N11503 0 diode
R11504 N11503 N11504 10
D11504 N11504 0 diode
R11505 N11504 N11505 10
D11505 N11505 0 diode
R11506 N11505 N11506 10
D11506 N11506 0 diode
R11507 N11506 N11507 10
D11507 N11507 0 diode
R11508 N11507 N11508 10
D11508 N11508 0 diode
R11509 N11508 N11509 10
D11509 N11509 0 diode
R11510 N11509 N11510 10
D11510 N11510 0 diode
R11511 N11510 N11511 10
D11511 N11511 0 diode
R11512 N11511 N11512 10
D11512 N11512 0 diode
R11513 N11512 N11513 10
D11513 N11513 0 diode
R11514 N11513 N11514 10
D11514 N11514 0 diode
R11515 N11514 N11515 10
D11515 N11515 0 diode
R11516 N11515 N11516 10
D11516 N11516 0 diode
R11517 N11516 N11517 10
D11517 N11517 0 diode
R11518 N11517 N11518 10
D11518 N11518 0 diode
R11519 N11518 N11519 10
D11519 N11519 0 diode
R11520 N11519 N11520 10
D11520 N11520 0 diode
R11521 N11520 N11521 10
D11521 N11521 0 diode
R11522 N11521 N11522 10
D11522 N11522 0 diode
R11523 N11522 N11523 10
D11523 N11523 0 diode
R11524 N11523 N11524 10
D11524 N11524 0 diode
R11525 N11524 N11525 10
D11525 N11525 0 diode
R11526 N11525 N11526 10
D11526 N11526 0 diode
R11527 N11526 N11527 10
D11527 N11527 0 diode
R11528 N11527 N11528 10
D11528 N11528 0 diode
R11529 N11528 N11529 10
D11529 N11529 0 diode
R11530 N11529 N11530 10
D11530 N11530 0 diode
R11531 N11530 N11531 10
D11531 N11531 0 diode
R11532 N11531 N11532 10
D11532 N11532 0 diode
R11533 N11532 N11533 10
D11533 N11533 0 diode
R11534 N11533 N11534 10
D11534 N11534 0 diode
R11535 N11534 N11535 10
D11535 N11535 0 diode
R11536 N11535 N11536 10
D11536 N11536 0 diode
R11537 N11536 N11537 10
D11537 N11537 0 diode
R11538 N11537 N11538 10
D11538 N11538 0 diode
R11539 N11538 N11539 10
D11539 N11539 0 diode
R11540 N11539 N11540 10
D11540 N11540 0 diode
R11541 N11540 N11541 10
D11541 N11541 0 diode
R11542 N11541 N11542 10
D11542 N11542 0 diode
R11543 N11542 N11543 10
D11543 N11543 0 diode
R11544 N11543 N11544 10
D11544 N11544 0 diode
R11545 N11544 N11545 10
D11545 N11545 0 diode
R11546 N11545 N11546 10
D11546 N11546 0 diode
R11547 N11546 N11547 10
D11547 N11547 0 diode
R11548 N11547 N11548 10
D11548 N11548 0 diode
R11549 N11548 N11549 10
D11549 N11549 0 diode
R11550 N11549 N11550 10
D11550 N11550 0 diode
R11551 N11550 N11551 10
D11551 N11551 0 diode
R11552 N11551 N11552 10
D11552 N11552 0 diode
R11553 N11552 N11553 10
D11553 N11553 0 diode
R11554 N11553 N11554 10
D11554 N11554 0 diode
R11555 N11554 N11555 10
D11555 N11555 0 diode
R11556 N11555 N11556 10
D11556 N11556 0 diode
R11557 N11556 N11557 10
D11557 N11557 0 diode
R11558 N11557 N11558 10
D11558 N11558 0 diode
R11559 N11558 N11559 10
D11559 N11559 0 diode
R11560 N11559 N11560 10
D11560 N11560 0 diode
R11561 N11560 N11561 10
D11561 N11561 0 diode
R11562 N11561 N11562 10
D11562 N11562 0 diode
R11563 N11562 N11563 10
D11563 N11563 0 diode
R11564 N11563 N11564 10
D11564 N11564 0 diode
R11565 N11564 N11565 10
D11565 N11565 0 diode
R11566 N11565 N11566 10
D11566 N11566 0 diode
R11567 N11566 N11567 10
D11567 N11567 0 diode
R11568 N11567 N11568 10
D11568 N11568 0 diode
R11569 N11568 N11569 10
D11569 N11569 0 diode
R11570 N11569 N11570 10
D11570 N11570 0 diode
R11571 N11570 N11571 10
D11571 N11571 0 diode
R11572 N11571 N11572 10
D11572 N11572 0 diode
R11573 N11572 N11573 10
D11573 N11573 0 diode
R11574 N11573 N11574 10
D11574 N11574 0 diode
R11575 N11574 N11575 10
D11575 N11575 0 diode
R11576 N11575 N11576 10
D11576 N11576 0 diode
R11577 N11576 N11577 10
D11577 N11577 0 diode
R11578 N11577 N11578 10
D11578 N11578 0 diode
R11579 N11578 N11579 10
D11579 N11579 0 diode
R11580 N11579 N11580 10
D11580 N11580 0 diode
R11581 N11580 N11581 10
D11581 N11581 0 diode
R11582 N11581 N11582 10
D11582 N11582 0 diode
R11583 N11582 N11583 10
D11583 N11583 0 diode
R11584 N11583 N11584 10
D11584 N11584 0 diode
R11585 N11584 N11585 10
D11585 N11585 0 diode
R11586 N11585 N11586 10
D11586 N11586 0 diode
R11587 N11586 N11587 10
D11587 N11587 0 diode
R11588 N11587 N11588 10
D11588 N11588 0 diode
R11589 N11588 N11589 10
D11589 N11589 0 diode
R11590 N11589 N11590 10
D11590 N11590 0 diode
R11591 N11590 N11591 10
D11591 N11591 0 diode
R11592 N11591 N11592 10
D11592 N11592 0 diode
R11593 N11592 N11593 10
D11593 N11593 0 diode
R11594 N11593 N11594 10
D11594 N11594 0 diode
R11595 N11594 N11595 10
D11595 N11595 0 diode
R11596 N11595 N11596 10
D11596 N11596 0 diode
R11597 N11596 N11597 10
D11597 N11597 0 diode
R11598 N11597 N11598 10
D11598 N11598 0 diode
R11599 N11598 N11599 10
D11599 N11599 0 diode
R11600 N11599 N11600 10
D11600 N11600 0 diode
R11601 N11600 N11601 10
D11601 N11601 0 diode
R11602 N11601 N11602 10
D11602 N11602 0 diode
R11603 N11602 N11603 10
D11603 N11603 0 diode
R11604 N11603 N11604 10
D11604 N11604 0 diode
R11605 N11604 N11605 10
D11605 N11605 0 diode
R11606 N11605 N11606 10
D11606 N11606 0 diode
R11607 N11606 N11607 10
D11607 N11607 0 diode
R11608 N11607 N11608 10
D11608 N11608 0 diode
R11609 N11608 N11609 10
D11609 N11609 0 diode
R11610 N11609 N11610 10
D11610 N11610 0 diode
R11611 N11610 N11611 10
D11611 N11611 0 diode
R11612 N11611 N11612 10
D11612 N11612 0 diode
R11613 N11612 N11613 10
D11613 N11613 0 diode
R11614 N11613 N11614 10
D11614 N11614 0 diode
R11615 N11614 N11615 10
D11615 N11615 0 diode
R11616 N11615 N11616 10
D11616 N11616 0 diode
R11617 N11616 N11617 10
D11617 N11617 0 diode
R11618 N11617 N11618 10
D11618 N11618 0 diode
R11619 N11618 N11619 10
D11619 N11619 0 diode
R11620 N11619 N11620 10
D11620 N11620 0 diode
R11621 N11620 N11621 10
D11621 N11621 0 diode
R11622 N11621 N11622 10
D11622 N11622 0 diode
R11623 N11622 N11623 10
D11623 N11623 0 diode
R11624 N11623 N11624 10
D11624 N11624 0 diode
R11625 N11624 N11625 10
D11625 N11625 0 diode
R11626 N11625 N11626 10
D11626 N11626 0 diode
R11627 N11626 N11627 10
D11627 N11627 0 diode
R11628 N11627 N11628 10
D11628 N11628 0 diode
R11629 N11628 N11629 10
D11629 N11629 0 diode
R11630 N11629 N11630 10
D11630 N11630 0 diode
R11631 N11630 N11631 10
D11631 N11631 0 diode
R11632 N11631 N11632 10
D11632 N11632 0 diode
R11633 N11632 N11633 10
D11633 N11633 0 diode
R11634 N11633 N11634 10
D11634 N11634 0 diode
R11635 N11634 N11635 10
D11635 N11635 0 diode
R11636 N11635 N11636 10
D11636 N11636 0 diode
R11637 N11636 N11637 10
D11637 N11637 0 diode
R11638 N11637 N11638 10
D11638 N11638 0 diode
R11639 N11638 N11639 10
D11639 N11639 0 diode
R11640 N11639 N11640 10
D11640 N11640 0 diode
R11641 N11640 N11641 10
D11641 N11641 0 diode
R11642 N11641 N11642 10
D11642 N11642 0 diode
R11643 N11642 N11643 10
D11643 N11643 0 diode
R11644 N11643 N11644 10
D11644 N11644 0 diode
R11645 N11644 N11645 10
D11645 N11645 0 diode
R11646 N11645 N11646 10
D11646 N11646 0 diode
R11647 N11646 N11647 10
D11647 N11647 0 diode
R11648 N11647 N11648 10
D11648 N11648 0 diode
R11649 N11648 N11649 10
D11649 N11649 0 diode
R11650 N11649 N11650 10
D11650 N11650 0 diode
R11651 N11650 N11651 10
D11651 N11651 0 diode
R11652 N11651 N11652 10
D11652 N11652 0 diode
R11653 N11652 N11653 10
D11653 N11653 0 diode
R11654 N11653 N11654 10
D11654 N11654 0 diode
R11655 N11654 N11655 10
D11655 N11655 0 diode
R11656 N11655 N11656 10
D11656 N11656 0 diode
R11657 N11656 N11657 10
D11657 N11657 0 diode
R11658 N11657 N11658 10
D11658 N11658 0 diode
R11659 N11658 N11659 10
D11659 N11659 0 diode
R11660 N11659 N11660 10
D11660 N11660 0 diode
R11661 N11660 N11661 10
D11661 N11661 0 diode
R11662 N11661 N11662 10
D11662 N11662 0 diode
R11663 N11662 N11663 10
D11663 N11663 0 diode
R11664 N11663 N11664 10
D11664 N11664 0 diode
R11665 N11664 N11665 10
D11665 N11665 0 diode
R11666 N11665 N11666 10
D11666 N11666 0 diode
R11667 N11666 N11667 10
D11667 N11667 0 diode
R11668 N11667 N11668 10
D11668 N11668 0 diode
R11669 N11668 N11669 10
D11669 N11669 0 diode
R11670 N11669 N11670 10
D11670 N11670 0 diode
R11671 N11670 N11671 10
D11671 N11671 0 diode
R11672 N11671 N11672 10
D11672 N11672 0 diode
R11673 N11672 N11673 10
D11673 N11673 0 diode
R11674 N11673 N11674 10
D11674 N11674 0 diode
R11675 N11674 N11675 10
D11675 N11675 0 diode
R11676 N11675 N11676 10
D11676 N11676 0 diode
R11677 N11676 N11677 10
D11677 N11677 0 diode
R11678 N11677 N11678 10
D11678 N11678 0 diode
R11679 N11678 N11679 10
D11679 N11679 0 diode
R11680 N11679 N11680 10
D11680 N11680 0 diode
R11681 N11680 N11681 10
D11681 N11681 0 diode
R11682 N11681 N11682 10
D11682 N11682 0 diode
R11683 N11682 N11683 10
D11683 N11683 0 diode
R11684 N11683 N11684 10
D11684 N11684 0 diode
R11685 N11684 N11685 10
D11685 N11685 0 diode
R11686 N11685 N11686 10
D11686 N11686 0 diode
R11687 N11686 N11687 10
D11687 N11687 0 diode
R11688 N11687 N11688 10
D11688 N11688 0 diode
R11689 N11688 N11689 10
D11689 N11689 0 diode
R11690 N11689 N11690 10
D11690 N11690 0 diode
R11691 N11690 N11691 10
D11691 N11691 0 diode
R11692 N11691 N11692 10
D11692 N11692 0 diode
R11693 N11692 N11693 10
D11693 N11693 0 diode
R11694 N11693 N11694 10
D11694 N11694 0 diode
R11695 N11694 N11695 10
D11695 N11695 0 diode
R11696 N11695 N11696 10
D11696 N11696 0 diode
R11697 N11696 N11697 10
D11697 N11697 0 diode
R11698 N11697 N11698 10
D11698 N11698 0 diode
R11699 N11698 N11699 10
D11699 N11699 0 diode
R11700 N11699 N11700 10
D11700 N11700 0 diode
R11701 N11700 N11701 10
D11701 N11701 0 diode
R11702 N11701 N11702 10
D11702 N11702 0 diode
R11703 N11702 N11703 10
D11703 N11703 0 diode
R11704 N11703 N11704 10
D11704 N11704 0 diode
R11705 N11704 N11705 10
D11705 N11705 0 diode
R11706 N11705 N11706 10
D11706 N11706 0 diode
R11707 N11706 N11707 10
D11707 N11707 0 diode
R11708 N11707 N11708 10
D11708 N11708 0 diode
R11709 N11708 N11709 10
D11709 N11709 0 diode
R11710 N11709 N11710 10
D11710 N11710 0 diode
R11711 N11710 N11711 10
D11711 N11711 0 diode
R11712 N11711 N11712 10
D11712 N11712 0 diode
R11713 N11712 N11713 10
D11713 N11713 0 diode
R11714 N11713 N11714 10
D11714 N11714 0 diode
R11715 N11714 N11715 10
D11715 N11715 0 diode
R11716 N11715 N11716 10
D11716 N11716 0 diode
R11717 N11716 N11717 10
D11717 N11717 0 diode
R11718 N11717 N11718 10
D11718 N11718 0 diode
R11719 N11718 N11719 10
D11719 N11719 0 diode
R11720 N11719 N11720 10
D11720 N11720 0 diode
R11721 N11720 N11721 10
D11721 N11721 0 diode
R11722 N11721 N11722 10
D11722 N11722 0 diode
R11723 N11722 N11723 10
D11723 N11723 0 diode
R11724 N11723 N11724 10
D11724 N11724 0 diode
R11725 N11724 N11725 10
D11725 N11725 0 diode
R11726 N11725 N11726 10
D11726 N11726 0 diode
R11727 N11726 N11727 10
D11727 N11727 0 diode
R11728 N11727 N11728 10
D11728 N11728 0 diode
R11729 N11728 N11729 10
D11729 N11729 0 diode
R11730 N11729 N11730 10
D11730 N11730 0 diode
R11731 N11730 N11731 10
D11731 N11731 0 diode
R11732 N11731 N11732 10
D11732 N11732 0 diode
R11733 N11732 N11733 10
D11733 N11733 0 diode
R11734 N11733 N11734 10
D11734 N11734 0 diode
R11735 N11734 N11735 10
D11735 N11735 0 diode
R11736 N11735 N11736 10
D11736 N11736 0 diode
R11737 N11736 N11737 10
D11737 N11737 0 diode
R11738 N11737 N11738 10
D11738 N11738 0 diode
R11739 N11738 N11739 10
D11739 N11739 0 diode
R11740 N11739 N11740 10
D11740 N11740 0 diode
R11741 N11740 N11741 10
D11741 N11741 0 diode
R11742 N11741 N11742 10
D11742 N11742 0 diode
R11743 N11742 N11743 10
D11743 N11743 0 diode
R11744 N11743 N11744 10
D11744 N11744 0 diode
R11745 N11744 N11745 10
D11745 N11745 0 diode
R11746 N11745 N11746 10
D11746 N11746 0 diode
R11747 N11746 N11747 10
D11747 N11747 0 diode
R11748 N11747 N11748 10
D11748 N11748 0 diode
R11749 N11748 N11749 10
D11749 N11749 0 diode
R11750 N11749 N11750 10
D11750 N11750 0 diode
R11751 N11750 N11751 10
D11751 N11751 0 diode
R11752 N11751 N11752 10
D11752 N11752 0 diode
R11753 N11752 N11753 10
D11753 N11753 0 diode
R11754 N11753 N11754 10
D11754 N11754 0 diode
R11755 N11754 N11755 10
D11755 N11755 0 diode
R11756 N11755 N11756 10
D11756 N11756 0 diode
R11757 N11756 N11757 10
D11757 N11757 0 diode
R11758 N11757 N11758 10
D11758 N11758 0 diode
R11759 N11758 N11759 10
D11759 N11759 0 diode
R11760 N11759 N11760 10
D11760 N11760 0 diode
R11761 N11760 N11761 10
D11761 N11761 0 diode
R11762 N11761 N11762 10
D11762 N11762 0 diode
R11763 N11762 N11763 10
D11763 N11763 0 diode
R11764 N11763 N11764 10
D11764 N11764 0 diode
R11765 N11764 N11765 10
D11765 N11765 0 diode
R11766 N11765 N11766 10
D11766 N11766 0 diode
R11767 N11766 N11767 10
D11767 N11767 0 diode
R11768 N11767 N11768 10
D11768 N11768 0 diode
R11769 N11768 N11769 10
D11769 N11769 0 diode
R11770 N11769 N11770 10
D11770 N11770 0 diode
R11771 N11770 N11771 10
D11771 N11771 0 diode
R11772 N11771 N11772 10
D11772 N11772 0 diode
R11773 N11772 N11773 10
D11773 N11773 0 diode
R11774 N11773 N11774 10
D11774 N11774 0 diode
R11775 N11774 N11775 10
D11775 N11775 0 diode
R11776 N11775 N11776 10
D11776 N11776 0 diode
R11777 N11776 N11777 10
D11777 N11777 0 diode
R11778 N11777 N11778 10
D11778 N11778 0 diode
R11779 N11778 N11779 10
D11779 N11779 0 diode
R11780 N11779 N11780 10
D11780 N11780 0 diode
R11781 N11780 N11781 10
D11781 N11781 0 diode
R11782 N11781 N11782 10
D11782 N11782 0 diode
R11783 N11782 N11783 10
D11783 N11783 0 diode
R11784 N11783 N11784 10
D11784 N11784 0 diode
R11785 N11784 N11785 10
D11785 N11785 0 diode
R11786 N11785 N11786 10
D11786 N11786 0 diode
R11787 N11786 N11787 10
D11787 N11787 0 diode
R11788 N11787 N11788 10
D11788 N11788 0 diode
R11789 N11788 N11789 10
D11789 N11789 0 diode
R11790 N11789 N11790 10
D11790 N11790 0 diode
R11791 N11790 N11791 10
D11791 N11791 0 diode
R11792 N11791 N11792 10
D11792 N11792 0 diode
R11793 N11792 N11793 10
D11793 N11793 0 diode
R11794 N11793 N11794 10
D11794 N11794 0 diode
R11795 N11794 N11795 10
D11795 N11795 0 diode
R11796 N11795 N11796 10
D11796 N11796 0 diode
R11797 N11796 N11797 10
D11797 N11797 0 diode
R11798 N11797 N11798 10
D11798 N11798 0 diode
R11799 N11798 N11799 10
D11799 N11799 0 diode
R11800 N11799 N11800 10
D11800 N11800 0 diode
R11801 N11800 N11801 10
D11801 N11801 0 diode
R11802 N11801 N11802 10
D11802 N11802 0 diode
R11803 N11802 N11803 10
D11803 N11803 0 diode
R11804 N11803 N11804 10
D11804 N11804 0 diode
R11805 N11804 N11805 10
D11805 N11805 0 diode
R11806 N11805 N11806 10
D11806 N11806 0 diode
R11807 N11806 N11807 10
D11807 N11807 0 diode
R11808 N11807 N11808 10
D11808 N11808 0 diode
R11809 N11808 N11809 10
D11809 N11809 0 diode
R11810 N11809 N11810 10
D11810 N11810 0 diode
R11811 N11810 N11811 10
D11811 N11811 0 diode
R11812 N11811 N11812 10
D11812 N11812 0 diode
R11813 N11812 N11813 10
D11813 N11813 0 diode
R11814 N11813 N11814 10
D11814 N11814 0 diode
R11815 N11814 N11815 10
D11815 N11815 0 diode
R11816 N11815 N11816 10
D11816 N11816 0 diode
R11817 N11816 N11817 10
D11817 N11817 0 diode
R11818 N11817 N11818 10
D11818 N11818 0 diode
R11819 N11818 N11819 10
D11819 N11819 0 diode
R11820 N11819 N11820 10
D11820 N11820 0 diode
R11821 N11820 N11821 10
D11821 N11821 0 diode
R11822 N11821 N11822 10
D11822 N11822 0 diode
R11823 N11822 N11823 10
D11823 N11823 0 diode
R11824 N11823 N11824 10
D11824 N11824 0 diode
R11825 N11824 N11825 10
D11825 N11825 0 diode
R11826 N11825 N11826 10
D11826 N11826 0 diode
R11827 N11826 N11827 10
D11827 N11827 0 diode
R11828 N11827 N11828 10
D11828 N11828 0 diode
R11829 N11828 N11829 10
D11829 N11829 0 diode
R11830 N11829 N11830 10
D11830 N11830 0 diode
R11831 N11830 N11831 10
D11831 N11831 0 diode
R11832 N11831 N11832 10
D11832 N11832 0 diode
R11833 N11832 N11833 10
D11833 N11833 0 diode
R11834 N11833 N11834 10
D11834 N11834 0 diode
R11835 N11834 N11835 10
D11835 N11835 0 diode
R11836 N11835 N11836 10
D11836 N11836 0 diode
R11837 N11836 N11837 10
D11837 N11837 0 diode
R11838 N11837 N11838 10
D11838 N11838 0 diode
R11839 N11838 N11839 10
D11839 N11839 0 diode
R11840 N11839 N11840 10
D11840 N11840 0 diode
R11841 N11840 N11841 10
D11841 N11841 0 diode
R11842 N11841 N11842 10
D11842 N11842 0 diode
R11843 N11842 N11843 10
D11843 N11843 0 diode
R11844 N11843 N11844 10
D11844 N11844 0 diode
R11845 N11844 N11845 10
D11845 N11845 0 diode
R11846 N11845 N11846 10
D11846 N11846 0 diode
R11847 N11846 N11847 10
D11847 N11847 0 diode
R11848 N11847 N11848 10
D11848 N11848 0 diode
R11849 N11848 N11849 10
D11849 N11849 0 diode
R11850 N11849 N11850 10
D11850 N11850 0 diode
R11851 N11850 N11851 10
D11851 N11851 0 diode
R11852 N11851 N11852 10
D11852 N11852 0 diode
R11853 N11852 N11853 10
D11853 N11853 0 diode
R11854 N11853 N11854 10
D11854 N11854 0 diode
R11855 N11854 N11855 10
D11855 N11855 0 diode
R11856 N11855 N11856 10
D11856 N11856 0 diode
R11857 N11856 N11857 10
D11857 N11857 0 diode
R11858 N11857 N11858 10
D11858 N11858 0 diode
R11859 N11858 N11859 10
D11859 N11859 0 diode
R11860 N11859 N11860 10
D11860 N11860 0 diode
R11861 N11860 N11861 10
D11861 N11861 0 diode
R11862 N11861 N11862 10
D11862 N11862 0 diode
R11863 N11862 N11863 10
D11863 N11863 0 diode
R11864 N11863 N11864 10
D11864 N11864 0 diode
R11865 N11864 N11865 10
D11865 N11865 0 diode
R11866 N11865 N11866 10
D11866 N11866 0 diode
R11867 N11866 N11867 10
D11867 N11867 0 diode
R11868 N11867 N11868 10
D11868 N11868 0 diode
R11869 N11868 N11869 10
D11869 N11869 0 diode
R11870 N11869 N11870 10
D11870 N11870 0 diode
R11871 N11870 N11871 10
D11871 N11871 0 diode
R11872 N11871 N11872 10
D11872 N11872 0 diode
R11873 N11872 N11873 10
D11873 N11873 0 diode
R11874 N11873 N11874 10
D11874 N11874 0 diode
R11875 N11874 N11875 10
D11875 N11875 0 diode
R11876 N11875 N11876 10
D11876 N11876 0 diode
R11877 N11876 N11877 10
D11877 N11877 0 diode
R11878 N11877 N11878 10
D11878 N11878 0 diode
R11879 N11878 N11879 10
D11879 N11879 0 diode
R11880 N11879 N11880 10
D11880 N11880 0 diode
R11881 N11880 N11881 10
D11881 N11881 0 diode
R11882 N11881 N11882 10
D11882 N11882 0 diode
R11883 N11882 N11883 10
D11883 N11883 0 diode
R11884 N11883 N11884 10
D11884 N11884 0 diode
R11885 N11884 N11885 10
D11885 N11885 0 diode
R11886 N11885 N11886 10
D11886 N11886 0 diode
R11887 N11886 N11887 10
D11887 N11887 0 diode
R11888 N11887 N11888 10
D11888 N11888 0 diode
R11889 N11888 N11889 10
D11889 N11889 0 diode
R11890 N11889 N11890 10
D11890 N11890 0 diode
R11891 N11890 N11891 10
D11891 N11891 0 diode
R11892 N11891 N11892 10
D11892 N11892 0 diode
R11893 N11892 N11893 10
D11893 N11893 0 diode
R11894 N11893 N11894 10
D11894 N11894 0 diode
R11895 N11894 N11895 10
D11895 N11895 0 diode
R11896 N11895 N11896 10
D11896 N11896 0 diode
R11897 N11896 N11897 10
D11897 N11897 0 diode
R11898 N11897 N11898 10
D11898 N11898 0 diode
R11899 N11898 N11899 10
D11899 N11899 0 diode
R11900 N11899 N11900 10
D11900 N11900 0 diode
R11901 N11900 N11901 10
D11901 N11901 0 diode
R11902 N11901 N11902 10
D11902 N11902 0 diode
R11903 N11902 N11903 10
D11903 N11903 0 diode
R11904 N11903 N11904 10
D11904 N11904 0 diode
R11905 N11904 N11905 10
D11905 N11905 0 diode
R11906 N11905 N11906 10
D11906 N11906 0 diode
R11907 N11906 N11907 10
D11907 N11907 0 diode
R11908 N11907 N11908 10
D11908 N11908 0 diode
R11909 N11908 N11909 10
D11909 N11909 0 diode
R11910 N11909 N11910 10
D11910 N11910 0 diode
R11911 N11910 N11911 10
D11911 N11911 0 diode
R11912 N11911 N11912 10
D11912 N11912 0 diode
R11913 N11912 N11913 10
D11913 N11913 0 diode
R11914 N11913 N11914 10
D11914 N11914 0 diode
R11915 N11914 N11915 10
D11915 N11915 0 diode
R11916 N11915 N11916 10
D11916 N11916 0 diode
R11917 N11916 N11917 10
D11917 N11917 0 diode
R11918 N11917 N11918 10
D11918 N11918 0 diode
R11919 N11918 N11919 10
D11919 N11919 0 diode
R11920 N11919 N11920 10
D11920 N11920 0 diode
R11921 N11920 N11921 10
D11921 N11921 0 diode
R11922 N11921 N11922 10
D11922 N11922 0 diode
R11923 N11922 N11923 10
D11923 N11923 0 diode
R11924 N11923 N11924 10
D11924 N11924 0 diode
R11925 N11924 N11925 10
D11925 N11925 0 diode
R11926 N11925 N11926 10
D11926 N11926 0 diode
R11927 N11926 N11927 10
D11927 N11927 0 diode
R11928 N11927 N11928 10
D11928 N11928 0 diode
R11929 N11928 N11929 10
D11929 N11929 0 diode
R11930 N11929 N11930 10
D11930 N11930 0 diode
R11931 N11930 N11931 10
D11931 N11931 0 diode
R11932 N11931 N11932 10
D11932 N11932 0 diode
R11933 N11932 N11933 10
D11933 N11933 0 diode
R11934 N11933 N11934 10
D11934 N11934 0 diode
R11935 N11934 N11935 10
D11935 N11935 0 diode
R11936 N11935 N11936 10
D11936 N11936 0 diode
R11937 N11936 N11937 10
D11937 N11937 0 diode
R11938 N11937 N11938 10
D11938 N11938 0 diode
R11939 N11938 N11939 10
D11939 N11939 0 diode
R11940 N11939 N11940 10
D11940 N11940 0 diode
R11941 N11940 N11941 10
D11941 N11941 0 diode
R11942 N11941 N11942 10
D11942 N11942 0 diode
R11943 N11942 N11943 10
D11943 N11943 0 diode
R11944 N11943 N11944 10
D11944 N11944 0 diode
R11945 N11944 N11945 10
D11945 N11945 0 diode
R11946 N11945 N11946 10
D11946 N11946 0 diode
R11947 N11946 N11947 10
D11947 N11947 0 diode
R11948 N11947 N11948 10
D11948 N11948 0 diode
R11949 N11948 N11949 10
D11949 N11949 0 diode
R11950 N11949 N11950 10
D11950 N11950 0 diode
R11951 N11950 N11951 10
D11951 N11951 0 diode
R11952 N11951 N11952 10
D11952 N11952 0 diode
R11953 N11952 N11953 10
D11953 N11953 0 diode
R11954 N11953 N11954 10
D11954 N11954 0 diode
R11955 N11954 N11955 10
D11955 N11955 0 diode
R11956 N11955 N11956 10
D11956 N11956 0 diode
R11957 N11956 N11957 10
D11957 N11957 0 diode
R11958 N11957 N11958 10
D11958 N11958 0 diode
R11959 N11958 N11959 10
D11959 N11959 0 diode
R11960 N11959 N11960 10
D11960 N11960 0 diode
R11961 N11960 N11961 10
D11961 N11961 0 diode
R11962 N11961 N11962 10
D11962 N11962 0 diode
R11963 N11962 N11963 10
D11963 N11963 0 diode
R11964 N11963 N11964 10
D11964 N11964 0 diode
R11965 N11964 N11965 10
D11965 N11965 0 diode
R11966 N11965 N11966 10
D11966 N11966 0 diode
R11967 N11966 N11967 10
D11967 N11967 0 diode
R11968 N11967 N11968 10
D11968 N11968 0 diode
R11969 N11968 N11969 10
D11969 N11969 0 diode
R11970 N11969 N11970 10
D11970 N11970 0 diode
R11971 N11970 N11971 10
D11971 N11971 0 diode
R11972 N11971 N11972 10
D11972 N11972 0 diode
R11973 N11972 N11973 10
D11973 N11973 0 diode
R11974 N11973 N11974 10
D11974 N11974 0 diode
R11975 N11974 N11975 10
D11975 N11975 0 diode
R11976 N11975 N11976 10
D11976 N11976 0 diode
R11977 N11976 N11977 10
D11977 N11977 0 diode
R11978 N11977 N11978 10
D11978 N11978 0 diode
R11979 N11978 N11979 10
D11979 N11979 0 diode
R11980 N11979 N11980 10
D11980 N11980 0 diode
R11981 N11980 N11981 10
D11981 N11981 0 diode
R11982 N11981 N11982 10
D11982 N11982 0 diode
R11983 N11982 N11983 10
D11983 N11983 0 diode
R11984 N11983 N11984 10
D11984 N11984 0 diode
R11985 N11984 N11985 10
D11985 N11985 0 diode
R11986 N11985 N11986 10
D11986 N11986 0 diode
R11987 N11986 N11987 10
D11987 N11987 0 diode
R11988 N11987 N11988 10
D11988 N11988 0 diode
R11989 N11988 N11989 10
D11989 N11989 0 diode
R11990 N11989 N11990 10
D11990 N11990 0 diode
R11991 N11990 N11991 10
D11991 N11991 0 diode
R11992 N11991 N11992 10
D11992 N11992 0 diode
R11993 N11992 N11993 10
D11993 N11993 0 diode
R11994 N11993 N11994 10
D11994 N11994 0 diode
R11995 N11994 N11995 10
D11995 N11995 0 diode
R11996 N11995 N11996 10
D11996 N11996 0 diode
R11997 N11996 N11997 10
D11997 N11997 0 diode
R11998 N11997 N11998 10
D11998 N11998 0 diode
R11999 N11998 N11999 10
D11999 N11999 0 diode
R12000 N11999 N12000 10
D12000 N12000 0 diode
R12001 N12000 N12001 10
D12001 N12001 0 diode
R12002 N12001 N12002 10
D12002 N12002 0 diode
R12003 N12002 N12003 10
D12003 N12003 0 diode
R12004 N12003 N12004 10
D12004 N12004 0 diode
R12005 N12004 N12005 10
D12005 N12005 0 diode
R12006 N12005 N12006 10
D12006 N12006 0 diode
R12007 N12006 N12007 10
D12007 N12007 0 diode
R12008 N12007 N12008 10
D12008 N12008 0 diode
R12009 N12008 N12009 10
D12009 N12009 0 diode
R12010 N12009 N12010 10
D12010 N12010 0 diode
R12011 N12010 N12011 10
D12011 N12011 0 diode
R12012 N12011 N12012 10
D12012 N12012 0 diode
R12013 N12012 N12013 10
D12013 N12013 0 diode
R12014 N12013 N12014 10
D12014 N12014 0 diode
R12015 N12014 N12015 10
D12015 N12015 0 diode
R12016 N12015 N12016 10
D12016 N12016 0 diode
R12017 N12016 N12017 10
D12017 N12017 0 diode
R12018 N12017 N12018 10
D12018 N12018 0 diode
R12019 N12018 N12019 10
D12019 N12019 0 diode
R12020 N12019 N12020 10
D12020 N12020 0 diode
R12021 N12020 N12021 10
D12021 N12021 0 diode
R12022 N12021 N12022 10
D12022 N12022 0 diode
R12023 N12022 N12023 10
D12023 N12023 0 diode
R12024 N12023 N12024 10
D12024 N12024 0 diode
R12025 N12024 N12025 10
D12025 N12025 0 diode
R12026 N12025 N12026 10
D12026 N12026 0 diode
R12027 N12026 N12027 10
D12027 N12027 0 diode
R12028 N12027 N12028 10
D12028 N12028 0 diode
R12029 N12028 N12029 10
D12029 N12029 0 diode
R12030 N12029 N12030 10
D12030 N12030 0 diode
R12031 N12030 N12031 10
D12031 N12031 0 diode
R12032 N12031 N12032 10
D12032 N12032 0 diode
R12033 N12032 N12033 10
D12033 N12033 0 diode
R12034 N12033 N12034 10
D12034 N12034 0 diode
R12035 N12034 N12035 10
D12035 N12035 0 diode
R12036 N12035 N12036 10
D12036 N12036 0 diode
R12037 N12036 N12037 10
D12037 N12037 0 diode
R12038 N12037 N12038 10
D12038 N12038 0 diode
R12039 N12038 N12039 10
D12039 N12039 0 diode
R12040 N12039 N12040 10
D12040 N12040 0 diode
R12041 N12040 N12041 10
D12041 N12041 0 diode
R12042 N12041 N12042 10
D12042 N12042 0 diode
R12043 N12042 N12043 10
D12043 N12043 0 diode
R12044 N12043 N12044 10
D12044 N12044 0 diode
R12045 N12044 N12045 10
D12045 N12045 0 diode
R12046 N12045 N12046 10
D12046 N12046 0 diode
R12047 N12046 N12047 10
D12047 N12047 0 diode
R12048 N12047 N12048 10
D12048 N12048 0 diode
R12049 N12048 N12049 10
D12049 N12049 0 diode
R12050 N12049 N12050 10
D12050 N12050 0 diode
R12051 N12050 N12051 10
D12051 N12051 0 diode
R12052 N12051 N12052 10
D12052 N12052 0 diode
R12053 N12052 N12053 10
D12053 N12053 0 diode
R12054 N12053 N12054 10
D12054 N12054 0 diode
R12055 N12054 N12055 10
D12055 N12055 0 diode
R12056 N12055 N12056 10
D12056 N12056 0 diode
R12057 N12056 N12057 10
D12057 N12057 0 diode
R12058 N12057 N12058 10
D12058 N12058 0 diode
R12059 N12058 N12059 10
D12059 N12059 0 diode
R12060 N12059 N12060 10
D12060 N12060 0 diode
R12061 N12060 N12061 10
D12061 N12061 0 diode
R12062 N12061 N12062 10
D12062 N12062 0 diode
R12063 N12062 N12063 10
D12063 N12063 0 diode
R12064 N12063 N12064 10
D12064 N12064 0 diode
R12065 N12064 N12065 10
D12065 N12065 0 diode
R12066 N12065 N12066 10
D12066 N12066 0 diode
R12067 N12066 N12067 10
D12067 N12067 0 diode
R12068 N12067 N12068 10
D12068 N12068 0 diode
R12069 N12068 N12069 10
D12069 N12069 0 diode
R12070 N12069 N12070 10
D12070 N12070 0 diode
R12071 N12070 N12071 10
D12071 N12071 0 diode
R12072 N12071 N12072 10
D12072 N12072 0 diode
R12073 N12072 N12073 10
D12073 N12073 0 diode
R12074 N12073 N12074 10
D12074 N12074 0 diode
R12075 N12074 N12075 10
D12075 N12075 0 diode
R12076 N12075 N12076 10
D12076 N12076 0 diode
R12077 N12076 N12077 10
D12077 N12077 0 diode
R12078 N12077 N12078 10
D12078 N12078 0 diode
R12079 N12078 N12079 10
D12079 N12079 0 diode
R12080 N12079 N12080 10
D12080 N12080 0 diode
R12081 N12080 N12081 10
D12081 N12081 0 diode
R12082 N12081 N12082 10
D12082 N12082 0 diode
R12083 N12082 N12083 10
D12083 N12083 0 diode
R12084 N12083 N12084 10
D12084 N12084 0 diode
R12085 N12084 N12085 10
D12085 N12085 0 diode
R12086 N12085 N12086 10
D12086 N12086 0 diode
R12087 N12086 N12087 10
D12087 N12087 0 diode
R12088 N12087 N12088 10
D12088 N12088 0 diode
R12089 N12088 N12089 10
D12089 N12089 0 diode
R12090 N12089 N12090 10
D12090 N12090 0 diode
R12091 N12090 N12091 10
D12091 N12091 0 diode
R12092 N12091 N12092 10
D12092 N12092 0 diode
R12093 N12092 N12093 10
D12093 N12093 0 diode
R12094 N12093 N12094 10
D12094 N12094 0 diode
R12095 N12094 N12095 10
D12095 N12095 0 diode
R12096 N12095 N12096 10
D12096 N12096 0 diode
R12097 N12096 N12097 10
D12097 N12097 0 diode
R12098 N12097 N12098 10
D12098 N12098 0 diode
R12099 N12098 N12099 10
D12099 N12099 0 diode
R12100 N12099 N12100 10
D12100 N12100 0 diode
R12101 N12100 N12101 10
D12101 N12101 0 diode
R12102 N12101 N12102 10
D12102 N12102 0 diode
R12103 N12102 N12103 10
D12103 N12103 0 diode
R12104 N12103 N12104 10
D12104 N12104 0 diode
R12105 N12104 N12105 10
D12105 N12105 0 diode
R12106 N12105 N12106 10
D12106 N12106 0 diode
R12107 N12106 N12107 10
D12107 N12107 0 diode
R12108 N12107 N12108 10
D12108 N12108 0 diode
R12109 N12108 N12109 10
D12109 N12109 0 diode
R12110 N12109 N12110 10
D12110 N12110 0 diode
R12111 N12110 N12111 10
D12111 N12111 0 diode
R12112 N12111 N12112 10
D12112 N12112 0 diode
R12113 N12112 N12113 10
D12113 N12113 0 diode
R12114 N12113 N12114 10
D12114 N12114 0 diode
R12115 N12114 N12115 10
D12115 N12115 0 diode
R12116 N12115 N12116 10
D12116 N12116 0 diode
R12117 N12116 N12117 10
D12117 N12117 0 diode
R12118 N12117 N12118 10
D12118 N12118 0 diode
R12119 N12118 N12119 10
D12119 N12119 0 diode
R12120 N12119 N12120 10
D12120 N12120 0 diode
R12121 N12120 N12121 10
D12121 N12121 0 diode
R12122 N12121 N12122 10
D12122 N12122 0 diode
R12123 N12122 N12123 10
D12123 N12123 0 diode
R12124 N12123 N12124 10
D12124 N12124 0 diode
R12125 N12124 N12125 10
D12125 N12125 0 diode
R12126 N12125 N12126 10
D12126 N12126 0 diode
R12127 N12126 N12127 10
D12127 N12127 0 diode
R12128 N12127 N12128 10
D12128 N12128 0 diode
R12129 N12128 N12129 10
D12129 N12129 0 diode
R12130 N12129 N12130 10
D12130 N12130 0 diode
R12131 N12130 N12131 10
D12131 N12131 0 diode
R12132 N12131 N12132 10
D12132 N12132 0 diode
R12133 N12132 N12133 10
D12133 N12133 0 diode
R12134 N12133 N12134 10
D12134 N12134 0 diode
R12135 N12134 N12135 10
D12135 N12135 0 diode
R12136 N12135 N12136 10
D12136 N12136 0 diode
R12137 N12136 N12137 10
D12137 N12137 0 diode
R12138 N12137 N12138 10
D12138 N12138 0 diode
R12139 N12138 N12139 10
D12139 N12139 0 diode
R12140 N12139 N12140 10
D12140 N12140 0 diode
R12141 N12140 N12141 10
D12141 N12141 0 diode
R12142 N12141 N12142 10
D12142 N12142 0 diode
R12143 N12142 N12143 10
D12143 N12143 0 diode
R12144 N12143 N12144 10
D12144 N12144 0 diode
R12145 N12144 N12145 10
D12145 N12145 0 diode
R12146 N12145 N12146 10
D12146 N12146 0 diode
R12147 N12146 N12147 10
D12147 N12147 0 diode
R12148 N12147 N12148 10
D12148 N12148 0 diode
R12149 N12148 N12149 10
D12149 N12149 0 diode
R12150 N12149 N12150 10
D12150 N12150 0 diode
R12151 N12150 N12151 10
D12151 N12151 0 diode
R12152 N12151 N12152 10
D12152 N12152 0 diode
R12153 N12152 N12153 10
D12153 N12153 0 diode
R12154 N12153 N12154 10
D12154 N12154 0 diode
R12155 N12154 N12155 10
D12155 N12155 0 diode
R12156 N12155 N12156 10
D12156 N12156 0 diode
R12157 N12156 N12157 10
D12157 N12157 0 diode
R12158 N12157 N12158 10
D12158 N12158 0 diode
R12159 N12158 N12159 10
D12159 N12159 0 diode
R12160 N12159 N12160 10
D12160 N12160 0 diode
R12161 N12160 N12161 10
D12161 N12161 0 diode
R12162 N12161 N12162 10
D12162 N12162 0 diode
R12163 N12162 N12163 10
D12163 N12163 0 diode
R12164 N12163 N12164 10
D12164 N12164 0 diode
R12165 N12164 N12165 10
D12165 N12165 0 diode
R12166 N12165 N12166 10
D12166 N12166 0 diode
R12167 N12166 N12167 10
D12167 N12167 0 diode
R12168 N12167 N12168 10
D12168 N12168 0 diode
R12169 N12168 N12169 10
D12169 N12169 0 diode
R12170 N12169 N12170 10
D12170 N12170 0 diode
R12171 N12170 N12171 10
D12171 N12171 0 diode
R12172 N12171 N12172 10
D12172 N12172 0 diode
R12173 N12172 N12173 10
D12173 N12173 0 diode
R12174 N12173 N12174 10
D12174 N12174 0 diode
R12175 N12174 N12175 10
D12175 N12175 0 diode
R12176 N12175 N12176 10
D12176 N12176 0 diode
R12177 N12176 N12177 10
D12177 N12177 0 diode
R12178 N12177 N12178 10
D12178 N12178 0 diode
R12179 N12178 N12179 10
D12179 N12179 0 diode
R12180 N12179 N12180 10
D12180 N12180 0 diode
R12181 N12180 N12181 10
D12181 N12181 0 diode
R12182 N12181 N12182 10
D12182 N12182 0 diode
R12183 N12182 N12183 10
D12183 N12183 0 diode
R12184 N12183 N12184 10
D12184 N12184 0 diode
R12185 N12184 N12185 10
D12185 N12185 0 diode
R12186 N12185 N12186 10
D12186 N12186 0 diode
R12187 N12186 N12187 10
D12187 N12187 0 diode
R12188 N12187 N12188 10
D12188 N12188 0 diode
R12189 N12188 N12189 10
D12189 N12189 0 diode
R12190 N12189 N12190 10
D12190 N12190 0 diode
R12191 N12190 N12191 10
D12191 N12191 0 diode
R12192 N12191 N12192 10
D12192 N12192 0 diode
R12193 N12192 N12193 10
D12193 N12193 0 diode
R12194 N12193 N12194 10
D12194 N12194 0 diode
R12195 N12194 N12195 10
D12195 N12195 0 diode
R12196 N12195 N12196 10
D12196 N12196 0 diode
R12197 N12196 N12197 10
D12197 N12197 0 diode
R12198 N12197 N12198 10
D12198 N12198 0 diode
R12199 N12198 N12199 10
D12199 N12199 0 diode
R12200 N12199 N12200 10
D12200 N12200 0 diode
R12201 N12200 N12201 10
D12201 N12201 0 diode
R12202 N12201 N12202 10
D12202 N12202 0 diode
R12203 N12202 N12203 10
D12203 N12203 0 diode
R12204 N12203 N12204 10
D12204 N12204 0 diode
R12205 N12204 N12205 10
D12205 N12205 0 diode
R12206 N12205 N12206 10
D12206 N12206 0 diode
R12207 N12206 N12207 10
D12207 N12207 0 diode
R12208 N12207 N12208 10
D12208 N12208 0 diode
R12209 N12208 N12209 10
D12209 N12209 0 diode
R12210 N12209 N12210 10
D12210 N12210 0 diode
R12211 N12210 N12211 10
D12211 N12211 0 diode
R12212 N12211 N12212 10
D12212 N12212 0 diode
R12213 N12212 N12213 10
D12213 N12213 0 diode
R12214 N12213 N12214 10
D12214 N12214 0 diode
R12215 N12214 N12215 10
D12215 N12215 0 diode
R12216 N12215 N12216 10
D12216 N12216 0 diode
R12217 N12216 N12217 10
D12217 N12217 0 diode
R12218 N12217 N12218 10
D12218 N12218 0 diode
R12219 N12218 N12219 10
D12219 N12219 0 diode
R12220 N12219 N12220 10
D12220 N12220 0 diode
R12221 N12220 N12221 10
D12221 N12221 0 diode
R12222 N12221 N12222 10
D12222 N12222 0 diode
R12223 N12222 N12223 10
D12223 N12223 0 diode
R12224 N12223 N12224 10
D12224 N12224 0 diode
R12225 N12224 N12225 10
D12225 N12225 0 diode
R12226 N12225 N12226 10
D12226 N12226 0 diode
R12227 N12226 N12227 10
D12227 N12227 0 diode
R12228 N12227 N12228 10
D12228 N12228 0 diode
R12229 N12228 N12229 10
D12229 N12229 0 diode
R12230 N12229 N12230 10
D12230 N12230 0 diode
R12231 N12230 N12231 10
D12231 N12231 0 diode
R12232 N12231 N12232 10
D12232 N12232 0 diode
R12233 N12232 N12233 10
D12233 N12233 0 diode
R12234 N12233 N12234 10
D12234 N12234 0 diode
R12235 N12234 N12235 10
D12235 N12235 0 diode
R12236 N12235 N12236 10
D12236 N12236 0 diode
R12237 N12236 N12237 10
D12237 N12237 0 diode
R12238 N12237 N12238 10
D12238 N12238 0 diode
R12239 N12238 N12239 10
D12239 N12239 0 diode
R12240 N12239 N12240 10
D12240 N12240 0 diode
R12241 N12240 N12241 10
D12241 N12241 0 diode
R12242 N12241 N12242 10
D12242 N12242 0 diode
R12243 N12242 N12243 10
D12243 N12243 0 diode
R12244 N12243 N12244 10
D12244 N12244 0 diode
R12245 N12244 N12245 10
D12245 N12245 0 diode
R12246 N12245 N12246 10
D12246 N12246 0 diode
R12247 N12246 N12247 10
D12247 N12247 0 diode
R12248 N12247 N12248 10
D12248 N12248 0 diode
R12249 N12248 N12249 10
D12249 N12249 0 diode
R12250 N12249 N12250 10
D12250 N12250 0 diode
R12251 N12250 N12251 10
D12251 N12251 0 diode
R12252 N12251 N12252 10
D12252 N12252 0 diode
R12253 N12252 N12253 10
D12253 N12253 0 diode
R12254 N12253 N12254 10
D12254 N12254 0 diode
R12255 N12254 N12255 10
D12255 N12255 0 diode
R12256 N12255 N12256 10
D12256 N12256 0 diode
R12257 N12256 N12257 10
D12257 N12257 0 diode
R12258 N12257 N12258 10
D12258 N12258 0 diode
R12259 N12258 N12259 10
D12259 N12259 0 diode
R12260 N12259 N12260 10
D12260 N12260 0 diode
R12261 N12260 N12261 10
D12261 N12261 0 diode
R12262 N12261 N12262 10
D12262 N12262 0 diode
R12263 N12262 N12263 10
D12263 N12263 0 diode
R12264 N12263 N12264 10
D12264 N12264 0 diode
R12265 N12264 N12265 10
D12265 N12265 0 diode
R12266 N12265 N12266 10
D12266 N12266 0 diode
R12267 N12266 N12267 10
D12267 N12267 0 diode
R12268 N12267 N12268 10
D12268 N12268 0 diode
R12269 N12268 N12269 10
D12269 N12269 0 diode
R12270 N12269 N12270 10
D12270 N12270 0 diode
R12271 N12270 N12271 10
D12271 N12271 0 diode
R12272 N12271 N12272 10
D12272 N12272 0 diode
R12273 N12272 N12273 10
D12273 N12273 0 diode
R12274 N12273 N12274 10
D12274 N12274 0 diode
R12275 N12274 N12275 10
D12275 N12275 0 diode
R12276 N12275 N12276 10
D12276 N12276 0 diode
R12277 N12276 N12277 10
D12277 N12277 0 diode
R12278 N12277 N12278 10
D12278 N12278 0 diode
R12279 N12278 N12279 10
D12279 N12279 0 diode
R12280 N12279 N12280 10
D12280 N12280 0 diode
R12281 N12280 N12281 10
D12281 N12281 0 diode
R12282 N12281 N12282 10
D12282 N12282 0 diode
R12283 N12282 N12283 10
D12283 N12283 0 diode
R12284 N12283 N12284 10
D12284 N12284 0 diode
R12285 N12284 N12285 10
D12285 N12285 0 diode
R12286 N12285 N12286 10
D12286 N12286 0 diode
R12287 N12286 N12287 10
D12287 N12287 0 diode
R12288 N12287 N12288 10
D12288 N12288 0 diode
R12289 N12288 N12289 10
D12289 N12289 0 diode
R12290 N12289 N12290 10
D12290 N12290 0 diode
R12291 N12290 N12291 10
D12291 N12291 0 diode
R12292 N12291 N12292 10
D12292 N12292 0 diode
R12293 N12292 N12293 10
D12293 N12293 0 diode
R12294 N12293 N12294 10
D12294 N12294 0 diode
R12295 N12294 N12295 10
D12295 N12295 0 diode
R12296 N12295 N12296 10
D12296 N12296 0 diode
R12297 N12296 N12297 10
D12297 N12297 0 diode
R12298 N12297 N12298 10
D12298 N12298 0 diode
R12299 N12298 N12299 10
D12299 N12299 0 diode
R12300 N12299 N12300 10
D12300 N12300 0 diode
R12301 N12300 N12301 10
D12301 N12301 0 diode
R12302 N12301 N12302 10
D12302 N12302 0 diode
R12303 N12302 N12303 10
D12303 N12303 0 diode
R12304 N12303 N12304 10
D12304 N12304 0 diode
R12305 N12304 N12305 10
D12305 N12305 0 diode
R12306 N12305 N12306 10
D12306 N12306 0 diode
R12307 N12306 N12307 10
D12307 N12307 0 diode
R12308 N12307 N12308 10
D12308 N12308 0 diode
R12309 N12308 N12309 10
D12309 N12309 0 diode
R12310 N12309 N12310 10
D12310 N12310 0 diode
R12311 N12310 N12311 10
D12311 N12311 0 diode
R12312 N12311 N12312 10
D12312 N12312 0 diode
R12313 N12312 N12313 10
D12313 N12313 0 diode
R12314 N12313 N12314 10
D12314 N12314 0 diode
R12315 N12314 N12315 10
D12315 N12315 0 diode
R12316 N12315 N12316 10
D12316 N12316 0 diode
R12317 N12316 N12317 10
D12317 N12317 0 diode
R12318 N12317 N12318 10
D12318 N12318 0 diode
R12319 N12318 N12319 10
D12319 N12319 0 diode
R12320 N12319 N12320 10
D12320 N12320 0 diode
R12321 N12320 N12321 10
D12321 N12321 0 diode
R12322 N12321 N12322 10
D12322 N12322 0 diode
R12323 N12322 N12323 10
D12323 N12323 0 diode
R12324 N12323 N12324 10
D12324 N12324 0 diode
R12325 N12324 N12325 10
D12325 N12325 0 diode
R12326 N12325 N12326 10
D12326 N12326 0 diode
R12327 N12326 N12327 10
D12327 N12327 0 diode
R12328 N12327 N12328 10
D12328 N12328 0 diode
R12329 N12328 N12329 10
D12329 N12329 0 diode
R12330 N12329 N12330 10
D12330 N12330 0 diode
R12331 N12330 N12331 10
D12331 N12331 0 diode
R12332 N12331 N12332 10
D12332 N12332 0 diode
R12333 N12332 N12333 10
D12333 N12333 0 diode
R12334 N12333 N12334 10
D12334 N12334 0 diode
R12335 N12334 N12335 10
D12335 N12335 0 diode
R12336 N12335 N12336 10
D12336 N12336 0 diode
R12337 N12336 N12337 10
D12337 N12337 0 diode
R12338 N12337 N12338 10
D12338 N12338 0 diode
R12339 N12338 N12339 10
D12339 N12339 0 diode
R12340 N12339 N12340 10
D12340 N12340 0 diode
R12341 N12340 N12341 10
D12341 N12341 0 diode
R12342 N12341 N12342 10
D12342 N12342 0 diode
R12343 N12342 N12343 10
D12343 N12343 0 diode
R12344 N12343 N12344 10
D12344 N12344 0 diode
R12345 N12344 N12345 10
D12345 N12345 0 diode
R12346 N12345 N12346 10
D12346 N12346 0 diode
R12347 N12346 N12347 10
D12347 N12347 0 diode
R12348 N12347 N12348 10
D12348 N12348 0 diode
R12349 N12348 N12349 10
D12349 N12349 0 diode
R12350 N12349 N12350 10
D12350 N12350 0 diode
R12351 N12350 N12351 10
D12351 N12351 0 diode
R12352 N12351 N12352 10
D12352 N12352 0 diode
R12353 N12352 N12353 10
D12353 N12353 0 diode
R12354 N12353 N12354 10
D12354 N12354 0 diode
R12355 N12354 N12355 10
D12355 N12355 0 diode
R12356 N12355 N12356 10
D12356 N12356 0 diode
R12357 N12356 N12357 10
D12357 N12357 0 diode
R12358 N12357 N12358 10
D12358 N12358 0 diode
R12359 N12358 N12359 10
D12359 N12359 0 diode
R12360 N12359 N12360 10
D12360 N12360 0 diode
R12361 N12360 N12361 10
D12361 N12361 0 diode
R12362 N12361 N12362 10
D12362 N12362 0 diode
R12363 N12362 N12363 10
D12363 N12363 0 diode
R12364 N12363 N12364 10
D12364 N12364 0 diode
R12365 N12364 N12365 10
D12365 N12365 0 diode
R12366 N12365 N12366 10
D12366 N12366 0 diode
R12367 N12366 N12367 10
D12367 N12367 0 diode
R12368 N12367 N12368 10
D12368 N12368 0 diode
R12369 N12368 N12369 10
D12369 N12369 0 diode
R12370 N12369 N12370 10
D12370 N12370 0 diode
R12371 N12370 N12371 10
D12371 N12371 0 diode
R12372 N12371 N12372 10
D12372 N12372 0 diode
R12373 N12372 N12373 10
D12373 N12373 0 diode
R12374 N12373 N12374 10
D12374 N12374 0 diode
R12375 N12374 N12375 10
D12375 N12375 0 diode
R12376 N12375 N12376 10
D12376 N12376 0 diode
R12377 N12376 N12377 10
D12377 N12377 0 diode
R12378 N12377 N12378 10
D12378 N12378 0 diode
R12379 N12378 N12379 10
D12379 N12379 0 diode
R12380 N12379 N12380 10
D12380 N12380 0 diode
R12381 N12380 N12381 10
D12381 N12381 0 diode
R12382 N12381 N12382 10
D12382 N12382 0 diode
R12383 N12382 N12383 10
D12383 N12383 0 diode
R12384 N12383 N12384 10
D12384 N12384 0 diode
R12385 N12384 N12385 10
D12385 N12385 0 diode
R12386 N12385 N12386 10
D12386 N12386 0 diode
R12387 N12386 N12387 10
D12387 N12387 0 diode
R12388 N12387 N12388 10
D12388 N12388 0 diode
R12389 N12388 N12389 10
D12389 N12389 0 diode
R12390 N12389 N12390 10
D12390 N12390 0 diode
R12391 N12390 N12391 10
D12391 N12391 0 diode
R12392 N12391 N12392 10
D12392 N12392 0 diode
R12393 N12392 N12393 10
D12393 N12393 0 diode
R12394 N12393 N12394 10
D12394 N12394 0 diode
R12395 N12394 N12395 10
D12395 N12395 0 diode
R12396 N12395 N12396 10
D12396 N12396 0 diode
R12397 N12396 N12397 10
D12397 N12397 0 diode
R12398 N12397 N12398 10
D12398 N12398 0 diode
R12399 N12398 N12399 10
D12399 N12399 0 diode
R12400 N12399 N12400 10
D12400 N12400 0 diode
R12401 N12400 N12401 10
D12401 N12401 0 diode
R12402 N12401 N12402 10
D12402 N12402 0 diode
R12403 N12402 N12403 10
D12403 N12403 0 diode
R12404 N12403 N12404 10
D12404 N12404 0 diode
R12405 N12404 N12405 10
D12405 N12405 0 diode
R12406 N12405 N12406 10
D12406 N12406 0 diode
R12407 N12406 N12407 10
D12407 N12407 0 diode
R12408 N12407 N12408 10
D12408 N12408 0 diode
R12409 N12408 N12409 10
D12409 N12409 0 diode
R12410 N12409 N12410 10
D12410 N12410 0 diode
R12411 N12410 N12411 10
D12411 N12411 0 diode
R12412 N12411 N12412 10
D12412 N12412 0 diode
R12413 N12412 N12413 10
D12413 N12413 0 diode
R12414 N12413 N12414 10
D12414 N12414 0 diode
R12415 N12414 N12415 10
D12415 N12415 0 diode
R12416 N12415 N12416 10
D12416 N12416 0 diode
R12417 N12416 N12417 10
D12417 N12417 0 diode
R12418 N12417 N12418 10
D12418 N12418 0 diode
R12419 N12418 N12419 10
D12419 N12419 0 diode
R12420 N12419 N12420 10
D12420 N12420 0 diode
R12421 N12420 N12421 10
D12421 N12421 0 diode
R12422 N12421 N12422 10
D12422 N12422 0 diode
R12423 N12422 N12423 10
D12423 N12423 0 diode
R12424 N12423 N12424 10
D12424 N12424 0 diode
R12425 N12424 N12425 10
D12425 N12425 0 diode
R12426 N12425 N12426 10
D12426 N12426 0 diode
R12427 N12426 N12427 10
D12427 N12427 0 diode
R12428 N12427 N12428 10
D12428 N12428 0 diode
R12429 N12428 N12429 10
D12429 N12429 0 diode
R12430 N12429 N12430 10
D12430 N12430 0 diode
R12431 N12430 N12431 10
D12431 N12431 0 diode
R12432 N12431 N12432 10
D12432 N12432 0 diode
R12433 N12432 N12433 10
D12433 N12433 0 diode
R12434 N12433 N12434 10
D12434 N12434 0 diode
R12435 N12434 N12435 10
D12435 N12435 0 diode
R12436 N12435 N12436 10
D12436 N12436 0 diode
R12437 N12436 N12437 10
D12437 N12437 0 diode
R12438 N12437 N12438 10
D12438 N12438 0 diode
R12439 N12438 N12439 10
D12439 N12439 0 diode
R12440 N12439 N12440 10
D12440 N12440 0 diode
R12441 N12440 N12441 10
D12441 N12441 0 diode
R12442 N12441 N12442 10
D12442 N12442 0 diode
R12443 N12442 N12443 10
D12443 N12443 0 diode
R12444 N12443 N12444 10
D12444 N12444 0 diode
R12445 N12444 N12445 10
D12445 N12445 0 diode
R12446 N12445 N12446 10
D12446 N12446 0 diode
R12447 N12446 N12447 10
D12447 N12447 0 diode
R12448 N12447 N12448 10
D12448 N12448 0 diode
R12449 N12448 N12449 10
D12449 N12449 0 diode
R12450 N12449 N12450 10
D12450 N12450 0 diode
R12451 N12450 N12451 10
D12451 N12451 0 diode
R12452 N12451 N12452 10
D12452 N12452 0 diode
R12453 N12452 N12453 10
D12453 N12453 0 diode
R12454 N12453 N12454 10
D12454 N12454 0 diode
R12455 N12454 N12455 10
D12455 N12455 0 diode
R12456 N12455 N12456 10
D12456 N12456 0 diode
R12457 N12456 N12457 10
D12457 N12457 0 diode
R12458 N12457 N12458 10
D12458 N12458 0 diode
R12459 N12458 N12459 10
D12459 N12459 0 diode
R12460 N12459 N12460 10
D12460 N12460 0 diode
R12461 N12460 N12461 10
D12461 N12461 0 diode
R12462 N12461 N12462 10
D12462 N12462 0 diode
R12463 N12462 N12463 10
D12463 N12463 0 diode
R12464 N12463 N12464 10
D12464 N12464 0 diode
R12465 N12464 N12465 10
D12465 N12465 0 diode
R12466 N12465 N12466 10
D12466 N12466 0 diode
R12467 N12466 N12467 10
D12467 N12467 0 diode
R12468 N12467 N12468 10
D12468 N12468 0 diode
R12469 N12468 N12469 10
D12469 N12469 0 diode
R12470 N12469 N12470 10
D12470 N12470 0 diode
R12471 N12470 N12471 10
D12471 N12471 0 diode
R12472 N12471 N12472 10
D12472 N12472 0 diode
R12473 N12472 N12473 10
D12473 N12473 0 diode
R12474 N12473 N12474 10
D12474 N12474 0 diode
R12475 N12474 N12475 10
D12475 N12475 0 diode
R12476 N12475 N12476 10
D12476 N12476 0 diode
R12477 N12476 N12477 10
D12477 N12477 0 diode
R12478 N12477 N12478 10
D12478 N12478 0 diode
R12479 N12478 N12479 10
D12479 N12479 0 diode
R12480 N12479 N12480 10
D12480 N12480 0 diode
R12481 N12480 N12481 10
D12481 N12481 0 diode
R12482 N12481 N12482 10
D12482 N12482 0 diode
R12483 N12482 N12483 10
D12483 N12483 0 diode
R12484 N12483 N12484 10
D12484 N12484 0 diode
R12485 N12484 N12485 10
D12485 N12485 0 diode
R12486 N12485 N12486 10
D12486 N12486 0 diode
R12487 N12486 N12487 10
D12487 N12487 0 diode
R12488 N12487 N12488 10
D12488 N12488 0 diode
R12489 N12488 N12489 10
D12489 N12489 0 diode
R12490 N12489 N12490 10
D12490 N12490 0 diode
R12491 N12490 N12491 10
D12491 N12491 0 diode
R12492 N12491 N12492 10
D12492 N12492 0 diode
R12493 N12492 N12493 10
D12493 N12493 0 diode
R12494 N12493 N12494 10
D12494 N12494 0 diode
R12495 N12494 N12495 10
D12495 N12495 0 diode
R12496 N12495 N12496 10
D12496 N12496 0 diode
R12497 N12496 N12497 10
D12497 N12497 0 diode
R12498 N12497 N12498 10
D12498 N12498 0 diode
R12499 N12498 N12499 10
D12499 N12499 0 diode
R12500 N12499 N12500 10
D12500 N12500 0 diode
R12501 N12500 N12501 10
D12501 N12501 0 diode
R12502 N12501 N12502 10
D12502 N12502 0 diode
R12503 N12502 N12503 10
D12503 N12503 0 diode
R12504 N12503 N12504 10
D12504 N12504 0 diode
R12505 N12504 N12505 10
D12505 N12505 0 diode
R12506 N12505 N12506 10
D12506 N12506 0 diode
R12507 N12506 N12507 10
D12507 N12507 0 diode
R12508 N12507 N12508 10
D12508 N12508 0 diode
R12509 N12508 N12509 10
D12509 N12509 0 diode
R12510 N12509 N12510 10
D12510 N12510 0 diode
R12511 N12510 N12511 10
D12511 N12511 0 diode
R12512 N12511 N12512 10
D12512 N12512 0 diode
R12513 N12512 N12513 10
D12513 N12513 0 diode
R12514 N12513 N12514 10
D12514 N12514 0 diode
R12515 N12514 N12515 10
D12515 N12515 0 diode
R12516 N12515 N12516 10
D12516 N12516 0 diode
R12517 N12516 N12517 10
D12517 N12517 0 diode
R12518 N12517 N12518 10
D12518 N12518 0 diode
R12519 N12518 N12519 10
D12519 N12519 0 diode
R12520 N12519 N12520 10
D12520 N12520 0 diode
R12521 N12520 N12521 10
D12521 N12521 0 diode
R12522 N12521 N12522 10
D12522 N12522 0 diode
R12523 N12522 N12523 10
D12523 N12523 0 diode
R12524 N12523 N12524 10
D12524 N12524 0 diode
R12525 N12524 N12525 10
D12525 N12525 0 diode
R12526 N12525 N12526 10
D12526 N12526 0 diode
R12527 N12526 N12527 10
D12527 N12527 0 diode
R12528 N12527 N12528 10
D12528 N12528 0 diode
R12529 N12528 N12529 10
D12529 N12529 0 diode
R12530 N12529 N12530 10
D12530 N12530 0 diode
R12531 N12530 N12531 10
D12531 N12531 0 diode
R12532 N12531 N12532 10
D12532 N12532 0 diode
R12533 N12532 N12533 10
D12533 N12533 0 diode
R12534 N12533 N12534 10
D12534 N12534 0 diode
R12535 N12534 N12535 10
D12535 N12535 0 diode
R12536 N12535 N12536 10
D12536 N12536 0 diode
R12537 N12536 N12537 10
D12537 N12537 0 diode
R12538 N12537 N12538 10
D12538 N12538 0 diode
R12539 N12538 N12539 10
D12539 N12539 0 diode
R12540 N12539 N12540 10
D12540 N12540 0 diode
R12541 N12540 N12541 10
D12541 N12541 0 diode
R12542 N12541 N12542 10
D12542 N12542 0 diode
R12543 N12542 N12543 10
D12543 N12543 0 diode
R12544 N12543 N12544 10
D12544 N12544 0 diode
R12545 N12544 N12545 10
D12545 N12545 0 diode
R12546 N12545 N12546 10
D12546 N12546 0 diode
R12547 N12546 N12547 10
D12547 N12547 0 diode
R12548 N12547 N12548 10
D12548 N12548 0 diode
R12549 N12548 N12549 10
D12549 N12549 0 diode
R12550 N12549 N12550 10
D12550 N12550 0 diode
R12551 N12550 N12551 10
D12551 N12551 0 diode
R12552 N12551 N12552 10
D12552 N12552 0 diode
R12553 N12552 N12553 10
D12553 N12553 0 diode
R12554 N12553 N12554 10
D12554 N12554 0 diode
R12555 N12554 N12555 10
D12555 N12555 0 diode
R12556 N12555 N12556 10
D12556 N12556 0 diode
R12557 N12556 N12557 10
D12557 N12557 0 diode
R12558 N12557 N12558 10
D12558 N12558 0 diode
R12559 N12558 N12559 10
D12559 N12559 0 diode
R12560 N12559 N12560 10
D12560 N12560 0 diode
R12561 N12560 N12561 10
D12561 N12561 0 diode
R12562 N12561 N12562 10
D12562 N12562 0 diode
R12563 N12562 N12563 10
D12563 N12563 0 diode
R12564 N12563 N12564 10
D12564 N12564 0 diode
R12565 N12564 N12565 10
D12565 N12565 0 diode
R12566 N12565 N12566 10
D12566 N12566 0 diode
R12567 N12566 N12567 10
D12567 N12567 0 diode
R12568 N12567 N12568 10
D12568 N12568 0 diode
R12569 N12568 N12569 10
D12569 N12569 0 diode
R12570 N12569 N12570 10
D12570 N12570 0 diode
R12571 N12570 N12571 10
D12571 N12571 0 diode
R12572 N12571 N12572 10
D12572 N12572 0 diode
R12573 N12572 N12573 10
D12573 N12573 0 diode
R12574 N12573 N12574 10
D12574 N12574 0 diode
R12575 N12574 N12575 10
D12575 N12575 0 diode
R12576 N12575 N12576 10
D12576 N12576 0 diode
R12577 N12576 N12577 10
D12577 N12577 0 diode
R12578 N12577 N12578 10
D12578 N12578 0 diode
R12579 N12578 N12579 10
D12579 N12579 0 diode
R12580 N12579 N12580 10
D12580 N12580 0 diode
R12581 N12580 N12581 10
D12581 N12581 0 diode
R12582 N12581 N12582 10
D12582 N12582 0 diode
R12583 N12582 N12583 10
D12583 N12583 0 diode
R12584 N12583 N12584 10
D12584 N12584 0 diode
R12585 N12584 N12585 10
D12585 N12585 0 diode
R12586 N12585 N12586 10
D12586 N12586 0 diode
R12587 N12586 N12587 10
D12587 N12587 0 diode
R12588 N12587 N12588 10
D12588 N12588 0 diode
R12589 N12588 N12589 10
D12589 N12589 0 diode
R12590 N12589 N12590 10
D12590 N12590 0 diode
R12591 N12590 N12591 10
D12591 N12591 0 diode
R12592 N12591 N12592 10
D12592 N12592 0 diode
R12593 N12592 N12593 10
D12593 N12593 0 diode
R12594 N12593 N12594 10
D12594 N12594 0 diode
R12595 N12594 N12595 10
D12595 N12595 0 diode
R12596 N12595 N12596 10
D12596 N12596 0 diode
R12597 N12596 N12597 10
D12597 N12597 0 diode
R12598 N12597 N12598 10
D12598 N12598 0 diode
R12599 N12598 N12599 10
D12599 N12599 0 diode
R12600 N12599 N12600 10
D12600 N12600 0 diode
R12601 N12600 N12601 10
D12601 N12601 0 diode
R12602 N12601 N12602 10
D12602 N12602 0 diode
R12603 N12602 N12603 10
D12603 N12603 0 diode
R12604 N12603 N12604 10
D12604 N12604 0 diode
R12605 N12604 N12605 10
D12605 N12605 0 diode
R12606 N12605 N12606 10
D12606 N12606 0 diode
R12607 N12606 N12607 10
D12607 N12607 0 diode
R12608 N12607 N12608 10
D12608 N12608 0 diode
R12609 N12608 N12609 10
D12609 N12609 0 diode
R12610 N12609 N12610 10
D12610 N12610 0 diode
R12611 N12610 N12611 10
D12611 N12611 0 diode
R12612 N12611 N12612 10
D12612 N12612 0 diode
R12613 N12612 N12613 10
D12613 N12613 0 diode
R12614 N12613 N12614 10
D12614 N12614 0 diode
R12615 N12614 N12615 10
D12615 N12615 0 diode
R12616 N12615 N12616 10
D12616 N12616 0 diode
R12617 N12616 N12617 10
D12617 N12617 0 diode
R12618 N12617 N12618 10
D12618 N12618 0 diode
R12619 N12618 N12619 10
D12619 N12619 0 diode
R12620 N12619 N12620 10
D12620 N12620 0 diode
R12621 N12620 N12621 10
D12621 N12621 0 diode
R12622 N12621 N12622 10
D12622 N12622 0 diode
R12623 N12622 N12623 10
D12623 N12623 0 diode
R12624 N12623 N12624 10
D12624 N12624 0 diode
R12625 N12624 N12625 10
D12625 N12625 0 diode
R12626 N12625 N12626 10
D12626 N12626 0 diode
R12627 N12626 N12627 10
D12627 N12627 0 diode
R12628 N12627 N12628 10
D12628 N12628 0 diode
R12629 N12628 N12629 10
D12629 N12629 0 diode
R12630 N12629 N12630 10
D12630 N12630 0 diode
R12631 N12630 N12631 10
D12631 N12631 0 diode
R12632 N12631 N12632 10
D12632 N12632 0 diode
R12633 N12632 N12633 10
D12633 N12633 0 diode
R12634 N12633 N12634 10
D12634 N12634 0 diode
R12635 N12634 N12635 10
D12635 N12635 0 diode
R12636 N12635 N12636 10
D12636 N12636 0 diode
R12637 N12636 N12637 10
D12637 N12637 0 diode
R12638 N12637 N12638 10
D12638 N12638 0 diode
R12639 N12638 N12639 10
D12639 N12639 0 diode
R12640 N12639 N12640 10
D12640 N12640 0 diode
R12641 N12640 N12641 10
D12641 N12641 0 diode
R12642 N12641 N12642 10
D12642 N12642 0 diode
R12643 N12642 N12643 10
D12643 N12643 0 diode
R12644 N12643 N12644 10
D12644 N12644 0 diode
R12645 N12644 N12645 10
D12645 N12645 0 diode
R12646 N12645 N12646 10
D12646 N12646 0 diode
R12647 N12646 N12647 10
D12647 N12647 0 diode
R12648 N12647 N12648 10
D12648 N12648 0 diode
R12649 N12648 N12649 10
D12649 N12649 0 diode
R12650 N12649 N12650 10
D12650 N12650 0 diode
R12651 N12650 N12651 10
D12651 N12651 0 diode
R12652 N12651 N12652 10
D12652 N12652 0 diode
R12653 N12652 N12653 10
D12653 N12653 0 diode
R12654 N12653 N12654 10
D12654 N12654 0 diode
R12655 N12654 N12655 10
D12655 N12655 0 diode
R12656 N12655 N12656 10
D12656 N12656 0 diode
R12657 N12656 N12657 10
D12657 N12657 0 diode
R12658 N12657 N12658 10
D12658 N12658 0 diode
R12659 N12658 N12659 10
D12659 N12659 0 diode
R12660 N12659 N12660 10
D12660 N12660 0 diode
R12661 N12660 N12661 10
D12661 N12661 0 diode
R12662 N12661 N12662 10
D12662 N12662 0 diode
R12663 N12662 N12663 10
D12663 N12663 0 diode
R12664 N12663 N12664 10
D12664 N12664 0 diode
R12665 N12664 N12665 10
D12665 N12665 0 diode
R12666 N12665 N12666 10
D12666 N12666 0 diode
R12667 N12666 N12667 10
D12667 N12667 0 diode
R12668 N12667 N12668 10
D12668 N12668 0 diode
R12669 N12668 N12669 10
D12669 N12669 0 diode
R12670 N12669 N12670 10
D12670 N12670 0 diode
R12671 N12670 N12671 10
D12671 N12671 0 diode
R12672 N12671 N12672 10
D12672 N12672 0 diode
R12673 N12672 N12673 10
D12673 N12673 0 diode
R12674 N12673 N12674 10
D12674 N12674 0 diode
R12675 N12674 N12675 10
D12675 N12675 0 diode
R12676 N12675 N12676 10
D12676 N12676 0 diode
R12677 N12676 N12677 10
D12677 N12677 0 diode
R12678 N12677 N12678 10
D12678 N12678 0 diode
R12679 N12678 N12679 10
D12679 N12679 0 diode
R12680 N12679 N12680 10
D12680 N12680 0 diode
R12681 N12680 N12681 10
D12681 N12681 0 diode
R12682 N12681 N12682 10
D12682 N12682 0 diode
R12683 N12682 N12683 10
D12683 N12683 0 diode
R12684 N12683 N12684 10
D12684 N12684 0 diode
R12685 N12684 N12685 10
D12685 N12685 0 diode
R12686 N12685 N12686 10
D12686 N12686 0 diode
R12687 N12686 N12687 10
D12687 N12687 0 diode
R12688 N12687 N12688 10
D12688 N12688 0 diode
R12689 N12688 N12689 10
D12689 N12689 0 diode
R12690 N12689 N12690 10
D12690 N12690 0 diode
R12691 N12690 N12691 10
D12691 N12691 0 diode
R12692 N12691 N12692 10
D12692 N12692 0 diode
R12693 N12692 N12693 10
D12693 N12693 0 diode
R12694 N12693 N12694 10
D12694 N12694 0 diode
R12695 N12694 N12695 10
D12695 N12695 0 diode
R12696 N12695 N12696 10
D12696 N12696 0 diode
R12697 N12696 N12697 10
D12697 N12697 0 diode
R12698 N12697 N12698 10
D12698 N12698 0 diode
R12699 N12698 N12699 10
D12699 N12699 0 diode
R12700 N12699 N12700 10
D12700 N12700 0 diode
R12701 N12700 N12701 10
D12701 N12701 0 diode
R12702 N12701 N12702 10
D12702 N12702 0 diode
R12703 N12702 N12703 10
D12703 N12703 0 diode
R12704 N12703 N12704 10
D12704 N12704 0 diode
R12705 N12704 N12705 10
D12705 N12705 0 diode
R12706 N12705 N12706 10
D12706 N12706 0 diode
R12707 N12706 N12707 10
D12707 N12707 0 diode
R12708 N12707 N12708 10
D12708 N12708 0 diode
R12709 N12708 N12709 10
D12709 N12709 0 diode
R12710 N12709 N12710 10
D12710 N12710 0 diode
R12711 N12710 N12711 10
D12711 N12711 0 diode
R12712 N12711 N12712 10
D12712 N12712 0 diode
R12713 N12712 N12713 10
D12713 N12713 0 diode
R12714 N12713 N12714 10
D12714 N12714 0 diode
R12715 N12714 N12715 10
D12715 N12715 0 diode
R12716 N12715 N12716 10
D12716 N12716 0 diode
R12717 N12716 N12717 10
D12717 N12717 0 diode
R12718 N12717 N12718 10
D12718 N12718 0 diode
R12719 N12718 N12719 10
D12719 N12719 0 diode
R12720 N12719 N12720 10
D12720 N12720 0 diode
R12721 N12720 N12721 10
D12721 N12721 0 diode
R12722 N12721 N12722 10
D12722 N12722 0 diode
R12723 N12722 N12723 10
D12723 N12723 0 diode
R12724 N12723 N12724 10
D12724 N12724 0 diode
R12725 N12724 N12725 10
D12725 N12725 0 diode
R12726 N12725 N12726 10
D12726 N12726 0 diode
R12727 N12726 N12727 10
D12727 N12727 0 diode
R12728 N12727 N12728 10
D12728 N12728 0 diode
R12729 N12728 N12729 10
D12729 N12729 0 diode
R12730 N12729 N12730 10
D12730 N12730 0 diode
R12731 N12730 N12731 10
D12731 N12731 0 diode
R12732 N12731 N12732 10
D12732 N12732 0 diode
R12733 N12732 N12733 10
D12733 N12733 0 diode
R12734 N12733 N12734 10
D12734 N12734 0 diode
R12735 N12734 N12735 10
D12735 N12735 0 diode
R12736 N12735 N12736 10
D12736 N12736 0 diode
R12737 N12736 N12737 10
D12737 N12737 0 diode
R12738 N12737 N12738 10
D12738 N12738 0 diode
R12739 N12738 N12739 10
D12739 N12739 0 diode
R12740 N12739 N12740 10
D12740 N12740 0 diode
R12741 N12740 N12741 10
D12741 N12741 0 diode
R12742 N12741 N12742 10
D12742 N12742 0 diode
R12743 N12742 N12743 10
D12743 N12743 0 diode
R12744 N12743 N12744 10
D12744 N12744 0 diode
R12745 N12744 N12745 10
D12745 N12745 0 diode
R12746 N12745 N12746 10
D12746 N12746 0 diode
R12747 N12746 N12747 10
D12747 N12747 0 diode
R12748 N12747 N12748 10
D12748 N12748 0 diode
R12749 N12748 N12749 10
D12749 N12749 0 diode
R12750 N12749 N12750 10
D12750 N12750 0 diode
R12751 N12750 N12751 10
D12751 N12751 0 diode
R12752 N12751 N12752 10
D12752 N12752 0 diode
R12753 N12752 N12753 10
D12753 N12753 0 diode
R12754 N12753 N12754 10
D12754 N12754 0 diode
R12755 N12754 N12755 10
D12755 N12755 0 diode
R12756 N12755 N12756 10
D12756 N12756 0 diode
R12757 N12756 N12757 10
D12757 N12757 0 diode
R12758 N12757 N12758 10
D12758 N12758 0 diode
R12759 N12758 N12759 10
D12759 N12759 0 diode
R12760 N12759 N12760 10
D12760 N12760 0 diode
R12761 N12760 N12761 10
D12761 N12761 0 diode
R12762 N12761 N12762 10
D12762 N12762 0 diode
R12763 N12762 N12763 10
D12763 N12763 0 diode
R12764 N12763 N12764 10
D12764 N12764 0 diode
R12765 N12764 N12765 10
D12765 N12765 0 diode
R12766 N12765 N12766 10
D12766 N12766 0 diode
R12767 N12766 N12767 10
D12767 N12767 0 diode
R12768 N12767 N12768 10
D12768 N12768 0 diode
R12769 N12768 N12769 10
D12769 N12769 0 diode
R12770 N12769 N12770 10
D12770 N12770 0 diode
R12771 N12770 N12771 10
D12771 N12771 0 diode
R12772 N12771 N12772 10
D12772 N12772 0 diode
R12773 N12772 N12773 10
D12773 N12773 0 diode
R12774 N12773 N12774 10
D12774 N12774 0 diode
R12775 N12774 N12775 10
D12775 N12775 0 diode
R12776 N12775 N12776 10
D12776 N12776 0 diode
R12777 N12776 N12777 10
D12777 N12777 0 diode
R12778 N12777 N12778 10
D12778 N12778 0 diode
R12779 N12778 N12779 10
D12779 N12779 0 diode
R12780 N12779 N12780 10
D12780 N12780 0 diode
R12781 N12780 N12781 10
D12781 N12781 0 diode
R12782 N12781 N12782 10
D12782 N12782 0 diode
R12783 N12782 N12783 10
D12783 N12783 0 diode
R12784 N12783 N12784 10
D12784 N12784 0 diode
R12785 N12784 N12785 10
D12785 N12785 0 diode
R12786 N12785 N12786 10
D12786 N12786 0 diode
R12787 N12786 N12787 10
D12787 N12787 0 diode
R12788 N12787 N12788 10
D12788 N12788 0 diode
R12789 N12788 N12789 10
D12789 N12789 0 diode
R12790 N12789 N12790 10
D12790 N12790 0 diode
R12791 N12790 N12791 10
D12791 N12791 0 diode
R12792 N12791 N12792 10
D12792 N12792 0 diode
R12793 N12792 N12793 10
D12793 N12793 0 diode
R12794 N12793 N12794 10
D12794 N12794 0 diode
R12795 N12794 N12795 10
D12795 N12795 0 diode
R12796 N12795 N12796 10
D12796 N12796 0 diode
R12797 N12796 N12797 10
D12797 N12797 0 diode
R12798 N12797 N12798 10
D12798 N12798 0 diode
R12799 N12798 N12799 10
D12799 N12799 0 diode
R12800 N12799 N12800 10
D12800 N12800 0 diode
R12801 N12800 N12801 10
D12801 N12801 0 diode
R12802 N12801 N12802 10
D12802 N12802 0 diode
R12803 N12802 N12803 10
D12803 N12803 0 diode
R12804 N12803 N12804 10
D12804 N12804 0 diode
R12805 N12804 N12805 10
D12805 N12805 0 diode
R12806 N12805 N12806 10
D12806 N12806 0 diode
R12807 N12806 N12807 10
D12807 N12807 0 diode
R12808 N12807 N12808 10
D12808 N12808 0 diode
R12809 N12808 N12809 10
D12809 N12809 0 diode
R12810 N12809 N12810 10
D12810 N12810 0 diode
R12811 N12810 N12811 10
D12811 N12811 0 diode
R12812 N12811 N12812 10
D12812 N12812 0 diode
R12813 N12812 N12813 10
D12813 N12813 0 diode
R12814 N12813 N12814 10
D12814 N12814 0 diode
R12815 N12814 N12815 10
D12815 N12815 0 diode
R12816 N12815 N12816 10
D12816 N12816 0 diode
R12817 N12816 N12817 10
D12817 N12817 0 diode
R12818 N12817 N12818 10
D12818 N12818 0 diode
R12819 N12818 N12819 10
D12819 N12819 0 diode
R12820 N12819 N12820 10
D12820 N12820 0 diode
R12821 N12820 N12821 10
D12821 N12821 0 diode
R12822 N12821 N12822 10
D12822 N12822 0 diode
R12823 N12822 N12823 10
D12823 N12823 0 diode
R12824 N12823 N12824 10
D12824 N12824 0 diode
R12825 N12824 N12825 10
D12825 N12825 0 diode
R12826 N12825 N12826 10
D12826 N12826 0 diode
R12827 N12826 N12827 10
D12827 N12827 0 diode
R12828 N12827 N12828 10
D12828 N12828 0 diode
R12829 N12828 N12829 10
D12829 N12829 0 diode
R12830 N12829 N12830 10
D12830 N12830 0 diode
R12831 N12830 N12831 10
D12831 N12831 0 diode
R12832 N12831 N12832 10
D12832 N12832 0 diode
R12833 N12832 N12833 10
D12833 N12833 0 diode
R12834 N12833 N12834 10
D12834 N12834 0 diode
R12835 N12834 N12835 10
D12835 N12835 0 diode
R12836 N12835 N12836 10
D12836 N12836 0 diode
R12837 N12836 N12837 10
D12837 N12837 0 diode
R12838 N12837 N12838 10
D12838 N12838 0 diode
R12839 N12838 N12839 10
D12839 N12839 0 diode
R12840 N12839 N12840 10
D12840 N12840 0 diode
R12841 N12840 N12841 10
D12841 N12841 0 diode
R12842 N12841 N12842 10
D12842 N12842 0 diode
R12843 N12842 N12843 10
D12843 N12843 0 diode
R12844 N12843 N12844 10
D12844 N12844 0 diode
R12845 N12844 N12845 10
D12845 N12845 0 diode
R12846 N12845 N12846 10
D12846 N12846 0 diode
R12847 N12846 N12847 10
D12847 N12847 0 diode
R12848 N12847 N12848 10
D12848 N12848 0 diode
R12849 N12848 N12849 10
D12849 N12849 0 diode
R12850 N12849 N12850 10
D12850 N12850 0 diode
R12851 N12850 N12851 10
D12851 N12851 0 diode
R12852 N12851 N12852 10
D12852 N12852 0 diode
R12853 N12852 N12853 10
D12853 N12853 0 diode
R12854 N12853 N12854 10
D12854 N12854 0 diode
R12855 N12854 N12855 10
D12855 N12855 0 diode
R12856 N12855 N12856 10
D12856 N12856 0 diode
R12857 N12856 N12857 10
D12857 N12857 0 diode
R12858 N12857 N12858 10
D12858 N12858 0 diode
R12859 N12858 N12859 10
D12859 N12859 0 diode
R12860 N12859 N12860 10
D12860 N12860 0 diode
R12861 N12860 N12861 10
D12861 N12861 0 diode
R12862 N12861 N12862 10
D12862 N12862 0 diode
R12863 N12862 N12863 10
D12863 N12863 0 diode
R12864 N12863 N12864 10
D12864 N12864 0 diode
R12865 N12864 N12865 10
D12865 N12865 0 diode
R12866 N12865 N12866 10
D12866 N12866 0 diode
R12867 N12866 N12867 10
D12867 N12867 0 diode
R12868 N12867 N12868 10
D12868 N12868 0 diode
R12869 N12868 N12869 10
D12869 N12869 0 diode
R12870 N12869 N12870 10
D12870 N12870 0 diode
R12871 N12870 N12871 10
D12871 N12871 0 diode
R12872 N12871 N12872 10
D12872 N12872 0 diode
R12873 N12872 N12873 10
D12873 N12873 0 diode
R12874 N12873 N12874 10
D12874 N12874 0 diode
R12875 N12874 N12875 10
D12875 N12875 0 diode
R12876 N12875 N12876 10
D12876 N12876 0 diode
R12877 N12876 N12877 10
D12877 N12877 0 diode
R12878 N12877 N12878 10
D12878 N12878 0 diode
R12879 N12878 N12879 10
D12879 N12879 0 diode
R12880 N12879 N12880 10
D12880 N12880 0 diode
R12881 N12880 N12881 10
D12881 N12881 0 diode
R12882 N12881 N12882 10
D12882 N12882 0 diode
R12883 N12882 N12883 10
D12883 N12883 0 diode
R12884 N12883 N12884 10
D12884 N12884 0 diode
R12885 N12884 N12885 10
D12885 N12885 0 diode
R12886 N12885 N12886 10
D12886 N12886 0 diode
R12887 N12886 N12887 10
D12887 N12887 0 diode
R12888 N12887 N12888 10
D12888 N12888 0 diode
R12889 N12888 N12889 10
D12889 N12889 0 diode
R12890 N12889 N12890 10
D12890 N12890 0 diode
R12891 N12890 N12891 10
D12891 N12891 0 diode
R12892 N12891 N12892 10
D12892 N12892 0 diode
R12893 N12892 N12893 10
D12893 N12893 0 diode
R12894 N12893 N12894 10
D12894 N12894 0 diode
R12895 N12894 N12895 10
D12895 N12895 0 diode
R12896 N12895 N12896 10
D12896 N12896 0 diode
R12897 N12896 N12897 10
D12897 N12897 0 diode
R12898 N12897 N12898 10
D12898 N12898 0 diode
R12899 N12898 N12899 10
D12899 N12899 0 diode
R12900 N12899 N12900 10
D12900 N12900 0 diode
R12901 N12900 N12901 10
D12901 N12901 0 diode
R12902 N12901 N12902 10
D12902 N12902 0 diode
R12903 N12902 N12903 10
D12903 N12903 0 diode
R12904 N12903 N12904 10
D12904 N12904 0 diode
R12905 N12904 N12905 10
D12905 N12905 0 diode
R12906 N12905 N12906 10
D12906 N12906 0 diode
R12907 N12906 N12907 10
D12907 N12907 0 diode
R12908 N12907 N12908 10
D12908 N12908 0 diode
R12909 N12908 N12909 10
D12909 N12909 0 diode
R12910 N12909 N12910 10
D12910 N12910 0 diode
R12911 N12910 N12911 10
D12911 N12911 0 diode
R12912 N12911 N12912 10
D12912 N12912 0 diode
R12913 N12912 N12913 10
D12913 N12913 0 diode
R12914 N12913 N12914 10
D12914 N12914 0 diode
R12915 N12914 N12915 10
D12915 N12915 0 diode
R12916 N12915 N12916 10
D12916 N12916 0 diode
R12917 N12916 N12917 10
D12917 N12917 0 diode
R12918 N12917 N12918 10
D12918 N12918 0 diode
R12919 N12918 N12919 10
D12919 N12919 0 diode
R12920 N12919 N12920 10
D12920 N12920 0 diode
R12921 N12920 N12921 10
D12921 N12921 0 diode
R12922 N12921 N12922 10
D12922 N12922 0 diode
R12923 N12922 N12923 10
D12923 N12923 0 diode
R12924 N12923 N12924 10
D12924 N12924 0 diode
R12925 N12924 N12925 10
D12925 N12925 0 diode
R12926 N12925 N12926 10
D12926 N12926 0 diode
R12927 N12926 N12927 10
D12927 N12927 0 diode
R12928 N12927 N12928 10
D12928 N12928 0 diode
R12929 N12928 N12929 10
D12929 N12929 0 diode
R12930 N12929 N12930 10
D12930 N12930 0 diode
R12931 N12930 N12931 10
D12931 N12931 0 diode
R12932 N12931 N12932 10
D12932 N12932 0 diode
R12933 N12932 N12933 10
D12933 N12933 0 diode
R12934 N12933 N12934 10
D12934 N12934 0 diode
R12935 N12934 N12935 10
D12935 N12935 0 diode
R12936 N12935 N12936 10
D12936 N12936 0 diode
R12937 N12936 N12937 10
D12937 N12937 0 diode
R12938 N12937 N12938 10
D12938 N12938 0 diode
R12939 N12938 N12939 10
D12939 N12939 0 diode
R12940 N12939 N12940 10
D12940 N12940 0 diode
R12941 N12940 N12941 10
D12941 N12941 0 diode
R12942 N12941 N12942 10
D12942 N12942 0 diode
R12943 N12942 N12943 10
D12943 N12943 0 diode
R12944 N12943 N12944 10
D12944 N12944 0 diode
R12945 N12944 N12945 10
D12945 N12945 0 diode
R12946 N12945 N12946 10
D12946 N12946 0 diode
R12947 N12946 N12947 10
D12947 N12947 0 diode
R12948 N12947 N12948 10
D12948 N12948 0 diode
R12949 N12948 N12949 10
D12949 N12949 0 diode
R12950 N12949 N12950 10
D12950 N12950 0 diode
R12951 N12950 N12951 10
D12951 N12951 0 diode
R12952 N12951 N12952 10
D12952 N12952 0 diode
R12953 N12952 N12953 10
D12953 N12953 0 diode
R12954 N12953 N12954 10
D12954 N12954 0 diode
R12955 N12954 N12955 10
D12955 N12955 0 diode
R12956 N12955 N12956 10
D12956 N12956 0 diode
R12957 N12956 N12957 10
D12957 N12957 0 diode
R12958 N12957 N12958 10
D12958 N12958 0 diode
R12959 N12958 N12959 10
D12959 N12959 0 diode
R12960 N12959 N12960 10
D12960 N12960 0 diode
R12961 N12960 N12961 10
D12961 N12961 0 diode
R12962 N12961 N12962 10
D12962 N12962 0 diode
R12963 N12962 N12963 10
D12963 N12963 0 diode
R12964 N12963 N12964 10
D12964 N12964 0 diode
R12965 N12964 N12965 10
D12965 N12965 0 diode
R12966 N12965 N12966 10
D12966 N12966 0 diode
R12967 N12966 N12967 10
D12967 N12967 0 diode
R12968 N12967 N12968 10
D12968 N12968 0 diode
R12969 N12968 N12969 10
D12969 N12969 0 diode
R12970 N12969 N12970 10
D12970 N12970 0 diode
R12971 N12970 N12971 10
D12971 N12971 0 diode
R12972 N12971 N12972 10
D12972 N12972 0 diode
R12973 N12972 N12973 10
D12973 N12973 0 diode
R12974 N12973 N12974 10
D12974 N12974 0 diode
R12975 N12974 N12975 10
D12975 N12975 0 diode
R12976 N12975 N12976 10
D12976 N12976 0 diode
R12977 N12976 N12977 10
D12977 N12977 0 diode
R12978 N12977 N12978 10
D12978 N12978 0 diode
R12979 N12978 N12979 10
D12979 N12979 0 diode
R12980 N12979 N12980 10
D12980 N12980 0 diode
R12981 N12980 N12981 10
D12981 N12981 0 diode
R12982 N12981 N12982 10
D12982 N12982 0 diode
R12983 N12982 N12983 10
D12983 N12983 0 diode
R12984 N12983 N12984 10
D12984 N12984 0 diode
R12985 N12984 N12985 10
D12985 N12985 0 diode
R12986 N12985 N12986 10
D12986 N12986 0 diode
R12987 N12986 N12987 10
D12987 N12987 0 diode
R12988 N12987 N12988 10
D12988 N12988 0 diode
R12989 N12988 N12989 10
D12989 N12989 0 diode
R12990 N12989 N12990 10
D12990 N12990 0 diode
R12991 N12990 N12991 10
D12991 N12991 0 diode
R12992 N12991 N12992 10
D12992 N12992 0 diode
R12993 N12992 N12993 10
D12993 N12993 0 diode
R12994 N12993 N12994 10
D12994 N12994 0 diode
R12995 N12994 N12995 10
D12995 N12995 0 diode
R12996 N12995 N12996 10
D12996 N12996 0 diode
R12997 N12996 N12997 10
D12997 N12997 0 diode
R12998 N12997 N12998 10
D12998 N12998 0 diode
R12999 N12998 N12999 10
D12999 N12999 0 diode
R13000 N12999 N13000 10
D13000 N13000 0 diode
R13001 N13000 N13001 10
D13001 N13001 0 diode
R13002 N13001 N13002 10
D13002 N13002 0 diode
R13003 N13002 N13003 10
D13003 N13003 0 diode
R13004 N13003 N13004 10
D13004 N13004 0 diode
R13005 N13004 N13005 10
D13005 N13005 0 diode
R13006 N13005 N13006 10
D13006 N13006 0 diode
R13007 N13006 N13007 10
D13007 N13007 0 diode
R13008 N13007 N13008 10
D13008 N13008 0 diode
R13009 N13008 N13009 10
D13009 N13009 0 diode
R13010 N13009 N13010 10
D13010 N13010 0 diode
R13011 N13010 N13011 10
D13011 N13011 0 diode
R13012 N13011 N13012 10
D13012 N13012 0 diode
R13013 N13012 N13013 10
D13013 N13013 0 diode
R13014 N13013 N13014 10
D13014 N13014 0 diode
R13015 N13014 N13015 10
D13015 N13015 0 diode
R13016 N13015 N13016 10
D13016 N13016 0 diode
R13017 N13016 N13017 10
D13017 N13017 0 diode
R13018 N13017 N13018 10
D13018 N13018 0 diode
R13019 N13018 N13019 10
D13019 N13019 0 diode
R13020 N13019 N13020 10
D13020 N13020 0 diode
R13021 N13020 N13021 10
D13021 N13021 0 diode
R13022 N13021 N13022 10
D13022 N13022 0 diode
R13023 N13022 N13023 10
D13023 N13023 0 diode
R13024 N13023 N13024 10
D13024 N13024 0 diode
R13025 N13024 N13025 10
D13025 N13025 0 diode
R13026 N13025 N13026 10
D13026 N13026 0 diode
R13027 N13026 N13027 10
D13027 N13027 0 diode
R13028 N13027 N13028 10
D13028 N13028 0 diode
R13029 N13028 N13029 10
D13029 N13029 0 diode
R13030 N13029 N13030 10
D13030 N13030 0 diode
R13031 N13030 N13031 10
D13031 N13031 0 diode
R13032 N13031 N13032 10
D13032 N13032 0 diode
R13033 N13032 N13033 10
D13033 N13033 0 diode
R13034 N13033 N13034 10
D13034 N13034 0 diode
R13035 N13034 N13035 10
D13035 N13035 0 diode
R13036 N13035 N13036 10
D13036 N13036 0 diode
R13037 N13036 N13037 10
D13037 N13037 0 diode
R13038 N13037 N13038 10
D13038 N13038 0 diode
R13039 N13038 N13039 10
D13039 N13039 0 diode
R13040 N13039 N13040 10
D13040 N13040 0 diode
R13041 N13040 N13041 10
D13041 N13041 0 diode
R13042 N13041 N13042 10
D13042 N13042 0 diode
R13043 N13042 N13043 10
D13043 N13043 0 diode
R13044 N13043 N13044 10
D13044 N13044 0 diode
R13045 N13044 N13045 10
D13045 N13045 0 diode
R13046 N13045 N13046 10
D13046 N13046 0 diode
R13047 N13046 N13047 10
D13047 N13047 0 diode
R13048 N13047 N13048 10
D13048 N13048 0 diode
R13049 N13048 N13049 10
D13049 N13049 0 diode
R13050 N13049 N13050 10
D13050 N13050 0 diode
R13051 N13050 N13051 10
D13051 N13051 0 diode
R13052 N13051 N13052 10
D13052 N13052 0 diode
R13053 N13052 N13053 10
D13053 N13053 0 diode
R13054 N13053 N13054 10
D13054 N13054 0 diode
R13055 N13054 N13055 10
D13055 N13055 0 diode
R13056 N13055 N13056 10
D13056 N13056 0 diode
R13057 N13056 N13057 10
D13057 N13057 0 diode
R13058 N13057 N13058 10
D13058 N13058 0 diode
R13059 N13058 N13059 10
D13059 N13059 0 diode
R13060 N13059 N13060 10
D13060 N13060 0 diode
R13061 N13060 N13061 10
D13061 N13061 0 diode
R13062 N13061 N13062 10
D13062 N13062 0 diode
R13063 N13062 N13063 10
D13063 N13063 0 diode
R13064 N13063 N13064 10
D13064 N13064 0 diode
R13065 N13064 N13065 10
D13065 N13065 0 diode
R13066 N13065 N13066 10
D13066 N13066 0 diode
R13067 N13066 N13067 10
D13067 N13067 0 diode
R13068 N13067 N13068 10
D13068 N13068 0 diode
R13069 N13068 N13069 10
D13069 N13069 0 diode
R13070 N13069 N13070 10
D13070 N13070 0 diode
R13071 N13070 N13071 10
D13071 N13071 0 diode
R13072 N13071 N13072 10
D13072 N13072 0 diode
R13073 N13072 N13073 10
D13073 N13073 0 diode
R13074 N13073 N13074 10
D13074 N13074 0 diode
R13075 N13074 N13075 10
D13075 N13075 0 diode
R13076 N13075 N13076 10
D13076 N13076 0 diode
R13077 N13076 N13077 10
D13077 N13077 0 diode
R13078 N13077 N13078 10
D13078 N13078 0 diode
R13079 N13078 N13079 10
D13079 N13079 0 diode
R13080 N13079 N13080 10
D13080 N13080 0 diode
R13081 N13080 N13081 10
D13081 N13081 0 diode
R13082 N13081 N13082 10
D13082 N13082 0 diode
R13083 N13082 N13083 10
D13083 N13083 0 diode
R13084 N13083 N13084 10
D13084 N13084 0 diode
R13085 N13084 N13085 10
D13085 N13085 0 diode
R13086 N13085 N13086 10
D13086 N13086 0 diode
R13087 N13086 N13087 10
D13087 N13087 0 diode
R13088 N13087 N13088 10
D13088 N13088 0 diode
R13089 N13088 N13089 10
D13089 N13089 0 diode
R13090 N13089 N13090 10
D13090 N13090 0 diode
R13091 N13090 N13091 10
D13091 N13091 0 diode
R13092 N13091 N13092 10
D13092 N13092 0 diode
R13093 N13092 N13093 10
D13093 N13093 0 diode
R13094 N13093 N13094 10
D13094 N13094 0 diode
R13095 N13094 N13095 10
D13095 N13095 0 diode
R13096 N13095 N13096 10
D13096 N13096 0 diode
R13097 N13096 N13097 10
D13097 N13097 0 diode
R13098 N13097 N13098 10
D13098 N13098 0 diode
R13099 N13098 N13099 10
D13099 N13099 0 diode
R13100 N13099 N13100 10
D13100 N13100 0 diode
R13101 N13100 N13101 10
D13101 N13101 0 diode
R13102 N13101 N13102 10
D13102 N13102 0 diode
R13103 N13102 N13103 10
D13103 N13103 0 diode
R13104 N13103 N13104 10
D13104 N13104 0 diode
R13105 N13104 N13105 10
D13105 N13105 0 diode
R13106 N13105 N13106 10
D13106 N13106 0 diode
R13107 N13106 N13107 10
D13107 N13107 0 diode
R13108 N13107 N13108 10
D13108 N13108 0 diode
R13109 N13108 N13109 10
D13109 N13109 0 diode
R13110 N13109 N13110 10
D13110 N13110 0 diode
R13111 N13110 N13111 10
D13111 N13111 0 diode
R13112 N13111 N13112 10
D13112 N13112 0 diode
R13113 N13112 N13113 10
D13113 N13113 0 diode
R13114 N13113 N13114 10
D13114 N13114 0 diode
R13115 N13114 N13115 10
D13115 N13115 0 diode
R13116 N13115 N13116 10
D13116 N13116 0 diode
R13117 N13116 N13117 10
D13117 N13117 0 diode
R13118 N13117 N13118 10
D13118 N13118 0 diode
R13119 N13118 N13119 10
D13119 N13119 0 diode
R13120 N13119 N13120 10
D13120 N13120 0 diode
R13121 N13120 N13121 10
D13121 N13121 0 diode
R13122 N13121 N13122 10
D13122 N13122 0 diode
R13123 N13122 N13123 10
D13123 N13123 0 diode
R13124 N13123 N13124 10
D13124 N13124 0 diode
R13125 N13124 N13125 10
D13125 N13125 0 diode
R13126 N13125 N13126 10
D13126 N13126 0 diode
R13127 N13126 N13127 10
D13127 N13127 0 diode
R13128 N13127 N13128 10
D13128 N13128 0 diode
R13129 N13128 N13129 10
D13129 N13129 0 diode
R13130 N13129 N13130 10
D13130 N13130 0 diode
R13131 N13130 N13131 10
D13131 N13131 0 diode
R13132 N13131 N13132 10
D13132 N13132 0 diode
R13133 N13132 N13133 10
D13133 N13133 0 diode
R13134 N13133 N13134 10
D13134 N13134 0 diode
R13135 N13134 N13135 10
D13135 N13135 0 diode
R13136 N13135 N13136 10
D13136 N13136 0 diode
R13137 N13136 N13137 10
D13137 N13137 0 diode
R13138 N13137 N13138 10
D13138 N13138 0 diode
R13139 N13138 N13139 10
D13139 N13139 0 diode
R13140 N13139 N13140 10
D13140 N13140 0 diode
R13141 N13140 N13141 10
D13141 N13141 0 diode
R13142 N13141 N13142 10
D13142 N13142 0 diode
R13143 N13142 N13143 10
D13143 N13143 0 diode
R13144 N13143 N13144 10
D13144 N13144 0 diode
R13145 N13144 N13145 10
D13145 N13145 0 diode
R13146 N13145 N13146 10
D13146 N13146 0 diode
R13147 N13146 N13147 10
D13147 N13147 0 diode
R13148 N13147 N13148 10
D13148 N13148 0 diode
R13149 N13148 N13149 10
D13149 N13149 0 diode
R13150 N13149 N13150 10
D13150 N13150 0 diode
R13151 N13150 N13151 10
D13151 N13151 0 diode
R13152 N13151 N13152 10
D13152 N13152 0 diode
R13153 N13152 N13153 10
D13153 N13153 0 diode
R13154 N13153 N13154 10
D13154 N13154 0 diode
R13155 N13154 N13155 10
D13155 N13155 0 diode
R13156 N13155 N13156 10
D13156 N13156 0 diode
R13157 N13156 N13157 10
D13157 N13157 0 diode
R13158 N13157 N13158 10
D13158 N13158 0 diode
R13159 N13158 N13159 10
D13159 N13159 0 diode
R13160 N13159 N13160 10
D13160 N13160 0 diode
R13161 N13160 N13161 10
D13161 N13161 0 diode
R13162 N13161 N13162 10
D13162 N13162 0 diode
R13163 N13162 N13163 10
D13163 N13163 0 diode
R13164 N13163 N13164 10
D13164 N13164 0 diode
R13165 N13164 N13165 10
D13165 N13165 0 diode
R13166 N13165 N13166 10
D13166 N13166 0 diode
R13167 N13166 N13167 10
D13167 N13167 0 diode
R13168 N13167 N13168 10
D13168 N13168 0 diode
R13169 N13168 N13169 10
D13169 N13169 0 diode
R13170 N13169 N13170 10
D13170 N13170 0 diode
R13171 N13170 N13171 10
D13171 N13171 0 diode
R13172 N13171 N13172 10
D13172 N13172 0 diode
R13173 N13172 N13173 10
D13173 N13173 0 diode
R13174 N13173 N13174 10
D13174 N13174 0 diode
R13175 N13174 N13175 10
D13175 N13175 0 diode
R13176 N13175 N13176 10
D13176 N13176 0 diode
R13177 N13176 N13177 10
D13177 N13177 0 diode
R13178 N13177 N13178 10
D13178 N13178 0 diode
R13179 N13178 N13179 10
D13179 N13179 0 diode
R13180 N13179 N13180 10
D13180 N13180 0 diode
R13181 N13180 N13181 10
D13181 N13181 0 diode
R13182 N13181 N13182 10
D13182 N13182 0 diode
R13183 N13182 N13183 10
D13183 N13183 0 diode
R13184 N13183 N13184 10
D13184 N13184 0 diode
R13185 N13184 N13185 10
D13185 N13185 0 diode
R13186 N13185 N13186 10
D13186 N13186 0 diode
R13187 N13186 N13187 10
D13187 N13187 0 diode
R13188 N13187 N13188 10
D13188 N13188 0 diode
R13189 N13188 N13189 10
D13189 N13189 0 diode
R13190 N13189 N13190 10
D13190 N13190 0 diode
R13191 N13190 N13191 10
D13191 N13191 0 diode
R13192 N13191 N13192 10
D13192 N13192 0 diode
R13193 N13192 N13193 10
D13193 N13193 0 diode
R13194 N13193 N13194 10
D13194 N13194 0 diode
R13195 N13194 N13195 10
D13195 N13195 0 diode
R13196 N13195 N13196 10
D13196 N13196 0 diode
R13197 N13196 N13197 10
D13197 N13197 0 diode
R13198 N13197 N13198 10
D13198 N13198 0 diode
R13199 N13198 N13199 10
D13199 N13199 0 diode
R13200 N13199 N13200 10
D13200 N13200 0 diode
R13201 N13200 N13201 10
D13201 N13201 0 diode
R13202 N13201 N13202 10
D13202 N13202 0 diode
R13203 N13202 N13203 10
D13203 N13203 0 diode
R13204 N13203 N13204 10
D13204 N13204 0 diode
R13205 N13204 N13205 10
D13205 N13205 0 diode
R13206 N13205 N13206 10
D13206 N13206 0 diode
R13207 N13206 N13207 10
D13207 N13207 0 diode
R13208 N13207 N13208 10
D13208 N13208 0 diode
R13209 N13208 N13209 10
D13209 N13209 0 diode
R13210 N13209 N13210 10
D13210 N13210 0 diode
R13211 N13210 N13211 10
D13211 N13211 0 diode
R13212 N13211 N13212 10
D13212 N13212 0 diode
R13213 N13212 N13213 10
D13213 N13213 0 diode
R13214 N13213 N13214 10
D13214 N13214 0 diode
R13215 N13214 N13215 10
D13215 N13215 0 diode
R13216 N13215 N13216 10
D13216 N13216 0 diode
R13217 N13216 N13217 10
D13217 N13217 0 diode
R13218 N13217 N13218 10
D13218 N13218 0 diode
R13219 N13218 N13219 10
D13219 N13219 0 diode
R13220 N13219 N13220 10
D13220 N13220 0 diode
R13221 N13220 N13221 10
D13221 N13221 0 diode
R13222 N13221 N13222 10
D13222 N13222 0 diode
R13223 N13222 N13223 10
D13223 N13223 0 diode
R13224 N13223 N13224 10
D13224 N13224 0 diode
R13225 N13224 N13225 10
D13225 N13225 0 diode
R13226 N13225 N13226 10
D13226 N13226 0 diode
R13227 N13226 N13227 10
D13227 N13227 0 diode
R13228 N13227 N13228 10
D13228 N13228 0 diode
R13229 N13228 N13229 10
D13229 N13229 0 diode
R13230 N13229 N13230 10
D13230 N13230 0 diode
R13231 N13230 N13231 10
D13231 N13231 0 diode
R13232 N13231 N13232 10
D13232 N13232 0 diode
R13233 N13232 N13233 10
D13233 N13233 0 diode
R13234 N13233 N13234 10
D13234 N13234 0 diode
R13235 N13234 N13235 10
D13235 N13235 0 diode
R13236 N13235 N13236 10
D13236 N13236 0 diode
R13237 N13236 N13237 10
D13237 N13237 0 diode
R13238 N13237 N13238 10
D13238 N13238 0 diode
R13239 N13238 N13239 10
D13239 N13239 0 diode
R13240 N13239 N13240 10
D13240 N13240 0 diode
R13241 N13240 N13241 10
D13241 N13241 0 diode
R13242 N13241 N13242 10
D13242 N13242 0 diode
R13243 N13242 N13243 10
D13243 N13243 0 diode
R13244 N13243 N13244 10
D13244 N13244 0 diode
R13245 N13244 N13245 10
D13245 N13245 0 diode
R13246 N13245 N13246 10
D13246 N13246 0 diode
R13247 N13246 N13247 10
D13247 N13247 0 diode
R13248 N13247 N13248 10
D13248 N13248 0 diode
R13249 N13248 N13249 10
D13249 N13249 0 diode
R13250 N13249 N13250 10
D13250 N13250 0 diode
R13251 N13250 N13251 10
D13251 N13251 0 diode
R13252 N13251 N13252 10
D13252 N13252 0 diode
R13253 N13252 N13253 10
D13253 N13253 0 diode
R13254 N13253 N13254 10
D13254 N13254 0 diode
R13255 N13254 N13255 10
D13255 N13255 0 diode
R13256 N13255 N13256 10
D13256 N13256 0 diode
R13257 N13256 N13257 10
D13257 N13257 0 diode
R13258 N13257 N13258 10
D13258 N13258 0 diode
R13259 N13258 N13259 10
D13259 N13259 0 diode
R13260 N13259 N13260 10
D13260 N13260 0 diode
R13261 N13260 N13261 10
D13261 N13261 0 diode
R13262 N13261 N13262 10
D13262 N13262 0 diode
R13263 N13262 N13263 10
D13263 N13263 0 diode
R13264 N13263 N13264 10
D13264 N13264 0 diode
R13265 N13264 N13265 10
D13265 N13265 0 diode
R13266 N13265 N13266 10
D13266 N13266 0 diode
R13267 N13266 N13267 10
D13267 N13267 0 diode
R13268 N13267 N13268 10
D13268 N13268 0 diode
R13269 N13268 N13269 10
D13269 N13269 0 diode
R13270 N13269 N13270 10
D13270 N13270 0 diode
R13271 N13270 N13271 10
D13271 N13271 0 diode
R13272 N13271 N13272 10
D13272 N13272 0 diode
R13273 N13272 N13273 10
D13273 N13273 0 diode
R13274 N13273 N13274 10
D13274 N13274 0 diode
R13275 N13274 N13275 10
D13275 N13275 0 diode
R13276 N13275 N13276 10
D13276 N13276 0 diode
R13277 N13276 N13277 10
D13277 N13277 0 diode
R13278 N13277 N13278 10
D13278 N13278 0 diode
R13279 N13278 N13279 10
D13279 N13279 0 diode
R13280 N13279 N13280 10
D13280 N13280 0 diode
R13281 N13280 N13281 10
D13281 N13281 0 diode
R13282 N13281 N13282 10
D13282 N13282 0 diode
R13283 N13282 N13283 10
D13283 N13283 0 diode
R13284 N13283 N13284 10
D13284 N13284 0 diode
R13285 N13284 N13285 10
D13285 N13285 0 diode
R13286 N13285 N13286 10
D13286 N13286 0 diode
R13287 N13286 N13287 10
D13287 N13287 0 diode
R13288 N13287 N13288 10
D13288 N13288 0 diode
R13289 N13288 N13289 10
D13289 N13289 0 diode
R13290 N13289 N13290 10
D13290 N13290 0 diode
R13291 N13290 N13291 10
D13291 N13291 0 diode
R13292 N13291 N13292 10
D13292 N13292 0 diode
R13293 N13292 N13293 10
D13293 N13293 0 diode
R13294 N13293 N13294 10
D13294 N13294 0 diode
R13295 N13294 N13295 10
D13295 N13295 0 diode
R13296 N13295 N13296 10
D13296 N13296 0 diode
R13297 N13296 N13297 10
D13297 N13297 0 diode
R13298 N13297 N13298 10
D13298 N13298 0 diode
R13299 N13298 N13299 10
D13299 N13299 0 diode
R13300 N13299 N13300 10
D13300 N13300 0 diode
R13301 N13300 N13301 10
D13301 N13301 0 diode
R13302 N13301 N13302 10
D13302 N13302 0 diode
R13303 N13302 N13303 10
D13303 N13303 0 diode
R13304 N13303 N13304 10
D13304 N13304 0 diode
R13305 N13304 N13305 10
D13305 N13305 0 diode
R13306 N13305 N13306 10
D13306 N13306 0 diode
R13307 N13306 N13307 10
D13307 N13307 0 diode
R13308 N13307 N13308 10
D13308 N13308 0 diode
R13309 N13308 N13309 10
D13309 N13309 0 diode
R13310 N13309 N13310 10
D13310 N13310 0 diode
R13311 N13310 N13311 10
D13311 N13311 0 diode
R13312 N13311 N13312 10
D13312 N13312 0 diode
R13313 N13312 N13313 10
D13313 N13313 0 diode
R13314 N13313 N13314 10
D13314 N13314 0 diode
R13315 N13314 N13315 10
D13315 N13315 0 diode
R13316 N13315 N13316 10
D13316 N13316 0 diode
R13317 N13316 N13317 10
D13317 N13317 0 diode
R13318 N13317 N13318 10
D13318 N13318 0 diode
R13319 N13318 N13319 10
D13319 N13319 0 diode
R13320 N13319 N13320 10
D13320 N13320 0 diode
R13321 N13320 N13321 10
D13321 N13321 0 diode
R13322 N13321 N13322 10
D13322 N13322 0 diode
R13323 N13322 N13323 10
D13323 N13323 0 diode
R13324 N13323 N13324 10
D13324 N13324 0 diode
R13325 N13324 N13325 10
D13325 N13325 0 diode
R13326 N13325 N13326 10
D13326 N13326 0 diode
R13327 N13326 N13327 10
D13327 N13327 0 diode
R13328 N13327 N13328 10
D13328 N13328 0 diode
R13329 N13328 N13329 10
D13329 N13329 0 diode
R13330 N13329 N13330 10
D13330 N13330 0 diode
R13331 N13330 N13331 10
D13331 N13331 0 diode
R13332 N13331 N13332 10
D13332 N13332 0 diode
R13333 N13332 N13333 10
D13333 N13333 0 diode
R13334 N13333 N13334 10
D13334 N13334 0 diode
R13335 N13334 N13335 10
D13335 N13335 0 diode
R13336 N13335 N13336 10
D13336 N13336 0 diode
R13337 N13336 N13337 10
D13337 N13337 0 diode
R13338 N13337 N13338 10
D13338 N13338 0 diode
R13339 N13338 N13339 10
D13339 N13339 0 diode
R13340 N13339 N13340 10
D13340 N13340 0 diode
R13341 N13340 N13341 10
D13341 N13341 0 diode
R13342 N13341 N13342 10
D13342 N13342 0 diode
R13343 N13342 N13343 10
D13343 N13343 0 diode
R13344 N13343 N13344 10
D13344 N13344 0 diode
R13345 N13344 N13345 10
D13345 N13345 0 diode
R13346 N13345 N13346 10
D13346 N13346 0 diode
R13347 N13346 N13347 10
D13347 N13347 0 diode
R13348 N13347 N13348 10
D13348 N13348 0 diode
R13349 N13348 N13349 10
D13349 N13349 0 diode
R13350 N13349 N13350 10
D13350 N13350 0 diode
R13351 N13350 N13351 10
D13351 N13351 0 diode
R13352 N13351 N13352 10
D13352 N13352 0 diode
R13353 N13352 N13353 10
D13353 N13353 0 diode
R13354 N13353 N13354 10
D13354 N13354 0 diode
R13355 N13354 N13355 10
D13355 N13355 0 diode
R13356 N13355 N13356 10
D13356 N13356 0 diode
R13357 N13356 N13357 10
D13357 N13357 0 diode
R13358 N13357 N13358 10
D13358 N13358 0 diode
R13359 N13358 N13359 10
D13359 N13359 0 diode
R13360 N13359 N13360 10
D13360 N13360 0 diode
R13361 N13360 N13361 10
D13361 N13361 0 diode
R13362 N13361 N13362 10
D13362 N13362 0 diode
R13363 N13362 N13363 10
D13363 N13363 0 diode
R13364 N13363 N13364 10
D13364 N13364 0 diode
R13365 N13364 N13365 10
D13365 N13365 0 diode
R13366 N13365 N13366 10
D13366 N13366 0 diode
R13367 N13366 N13367 10
D13367 N13367 0 diode
R13368 N13367 N13368 10
D13368 N13368 0 diode
R13369 N13368 N13369 10
D13369 N13369 0 diode
R13370 N13369 N13370 10
D13370 N13370 0 diode
R13371 N13370 N13371 10
D13371 N13371 0 diode
R13372 N13371 N13372 10
D13372 N13372 0 diode
R13373 N13372 N13373 10
D13373 N13373 0 diode
R13374 N13373 N13374 10
D13374 N13374 0 diode
R13375 N13374 N13375 10
D13375 N13375 0 diode
R13376 N13375 N13376 10
D13376 N13376 0 diode
R13377 N13376 N13377 10
D13377 N13377 0 diode
R13378 N13377 N13378 10
D13378 N13378 0 diode
R13379 N13378 N13379 10
D13379 N13379 0 diode
R13380 N13379 N13380 10
D13380 N13380 0 diode
R13381 N13380 N13381 10
D13381 N13381 0 diode
R13382 N13381 N13382 10
D13382 N13382 0 diode
R13383 N13382 N13383 10
D13383 N13383 0 diode
R13384 N13383 N13384 10
D13384 N13384 0 diode
R13385 N13384 N13385 10
D13385 N13385 0 diode
R13386 N13385 N13386 10
D13386 N13386 0 diode
R13387 N13386 N13387 10
D13387 N13387 0 diode
R13388 N13387 N13388 10
D13388 N13388 0 diode
R13389 N13388 N13389 10
D13389 N13389 0 diode
R13390 N13389 N13390 10
D13390 N13390 0 diode
R13391 N13390 N13391 10
D13391 N13391 0 diode
R13392 N13391 N13392 10
D13392 N13392 0 diode
R13393 N13392 N13393 10
D13393 N13393 0 diode
R13394 N13393 N13394 10
D13394 N13394 0 diode
R13395 N13394 N13395 10
D13395 N13395 0 diode
R13396 N13395 N13396 10
D13396 N13396 0 diode
R13397 N13396 N13397 10
D13397 N13397 0 diode
R13398 N13397 N13398 10
D13398 N13398 0 diode
R13399 N13398 N13399 10
D13399 N13399 0 diode
R13400 N13399 N13400 10
D13400 N13400 0 diode
R13401 N13400 N13401 10
D13401 N13401 0 diode
R13402 N13401 N13402 10
D13402 N13402 0 diode
R13403 N13402 N13403 10
D13403 N13403 0 diode
R13404 N13403 N13404 10
D13404 N13404 0 diode
R13405 N13404 N13405 10
D13405 N13405 0 diode
R13406 N13405 N13406 10
D13406 N13406 0 diode
R13407 N13406 N13407 10
D13407 N13407 0 diode
R13408 N13407 N13408 10
D13408 N13408 0 diode
R13409 N13408 N13409 10
D13409 N13409 0 diode
R13410 N13409 N13410 10
D13410 N13410 0 diode
R13411 N13410 N13411 10
D13411 N13411 0 diode
R13412 N13411 N13412 10
D13412 N13412 0 diode
R13413 N13412 N13413 10
D13413 N13413 0 diode
R13414 N13413 N13414 10
D13414 N13414 0 diode
R13415 N13414 N13415 10
D13415 N13415 0 diode
R13416 N13415 N13416 10
D13416 N13416 0 diode
R13417 N13416 N13417 10
D13417 N13417 0 diode
R13418 N13417 N13418 10
D13418 N13418 0 diode
R13419 N13418 N13419 10
D13419 N13419 0 diode
R13420 N13419 N13420 10
D13420 N13420 0 diode
R13421 N13420 N13421 10
D13421 N13421 0 diode
R13422 N13421 N13422 10
D13422 N13422 0 diode
R13423 N13422 N13423 10
D13423 N13423 0 diode
R13424 N13423 N13424 10
D13424 N13424 0 diode
R13425 N13424 N13425 10
D13425 N13425 0 diode
R13426 N13425 N13426 10
D13426 N13426 0 diode
R13427 N13426 N13427 10
D13427 N13427 0 diode
R13428 N13427 N13428 10
D13428 N13428 0 diode
R13429 N13428 N13429 10
D13429 N13429 0 diode
R13430 N13429 N13430 10
D13430 N13430 0 diode
R13431 N13430 N13431 10
D13431 N13431 0 diode
R13432 N13431 N13432 10
D13432 N13432 0 diode
R13433 N13432 N13433 10
D13433 N13433 0 diode
R13434 N13433 N13434 10
D13434 N13434 0 diode
R13435 N13434 N13435 10
D13435 N13435 0 diode
R13436 N13435 N13436 10
D13436 N13436 0 diode
R13437 N13436 N13437 10
D13437 N13437 0 diode
R13438 N13437 N13438 10
D13438 N13438 0 diode
R13439 N13438 N13439 10
D13439 N13439 0 diode
R13440 N13439 N13440 10
D13440 N13440 0 diode
R13441 N13440 N13441 10
D13441 N13441 0 diode
R13442 N13441 N13442 10
D13442 N13442 0 diode
R13443 N13442 N13443 10
D13443 N13443 0 diode
R13444 N13443 N13444 10
D13444 N13444 0 diode
R13445 N13444 N13445 10
D13445 N13445 0 diode
R13446 N13445 N13446 10
D13446 N13446 0 diode
R13447 N13446 N13447 10
D13447 N13447 0 diode
R13448 N13447 N13448 10
D13448 N13448 0 diode
R13449 N13448 N13449 10
D13449 N13449 0 diode
R13450 N13449 N13450 10
D13450 N13450 0 diode
R13451 N13450 N13451 10
D13451 N13451 0 diode
R13452 N13451 N13452 10
D13452 N13452 0 diode
R13453 N13452 N13453 10
D13453 N13453 0 diode
R13454 N13453 N13454 10
D13454 N13454 0 diode
R13455 N13454 N13455 10
D13455 N13455 0 diode
R13456 N13455 N13456 10
D13456 N13456 0 diode
R13457 N13456 N13457 10
D13457 N13457 0 diode
R13458 N13457 N13458 10
D13458 N13458 0 diode
R13459 N13458 N13459 10
D13459 N13459 0 diode
R13460 N13459 N13460 10
D13460 N13460 0 diode
R13461 N13460 N13461 10
D13461 N13461 0 diode
R13462 N13461 N13462 10
D13462 N13462 0 diode
R13463 N13462 N13463 10
D13463 N13463 0 diode
R13464 N13463 N13464 10
D13464 N13464 0 diode
R13465 N13464 N13465 10
D13465 N13465 0 diode
R13466 N13465 N13466 10
D13466 N13466 0 diode
R13467 N13466 N13467 10
D13467 N13467 0 diode
R13468 N13467 N13468 10
D13468 N13468 0 diode
R13469 N13468 N13469 10
D13469 N13469 0 diode
R13470 N13469 N13470 10
D13470 N13470 0 diode
R13471 N13470 N13471 10
D13471 N13471 0 diode
R13472 N13471 N13472 10
D13472 N13472 0 diode
R13473 N13472 N13473 10
D13473 N13473 0 diode
R13474 N13473 N13474 10
D13474 N13474 0 diode
R13475 N13474 N13475 10
D13475 N13475 0 diode
R13476 N13475 N13476 10
D13476 N13476 0 diode
R13477 N13476 N13477 10
D13477 N13477 0 diode
R13478 N13477 N13478 10
D13478 N13478 0 diode
R13479 N13478 N13479 10
D13479 N13479 0 diode
R13480 N13479 N13480 10
D13480 N13480 0 diode
R13481 N13480 N13481 10
D13481 N13481 0 diode
R13482 N13481 N13482 10
D13482 N13482 0 diode
R13483 N13482 N13483 10
D13483 N13483 0 diode
R13484 N13483 N13484 10
D13484 N13484 0 diode
R13485 N13484 N13485 10
D13485 N13485 0 diode
R13486 N13485 N13486 10
D13486 N13486 0 diode
R13487 N13486 N13487 10
D13487 N13487 0 diode
R13488 N13487 N13488 10
D13488 N13488 0 diode
R13489 N13488 N13489 10
D13489 N13489 0 diode
R13490 N13489 N13490 10
D13490 N13490 0 diode
R13491 N13490 N13491 10
D13491 N13491 0 diode
R13492 N13491 N13492 10
D13492 N13492 0 diode
R13493 N13492 N13493 10
D13493 N13493 0 diode
R13494 N13493 N13494 10
D13494 N13494 0 diode
R13495 N13494 N13495 10
D13495 N13495 0 diode
R13496 N13495 N13496 10
D13496 N13496 0 diode
R13497 N13496 N13497 10
D13497 N13497 0 diode
R13498 N13497 N13498 10
D13498 N13498 0 diode
R13499 N13498 N13499 10
D13499 N13499 0 diode
R13500 N13499 N13500 10
D13500 N13500 0 diode
R13501 N13500 N13501 10
D13501 N13501 0 diode
R13502 N13501 N13502 10
D13502 N13502 0 diode
R13503 N13502 N13503 10
D13503 N13503 0 diode
R13504 N13503 N13504 10
D13504 N13504 0 diode
R13505 N13504 N13505 10
D13505 N13505 0 diode
R13506 N13505 N13506 10
D13506 N13506 0 diode
R13507 N13506 N13507 10
D13507 N13507 0 diode
R13508 N13507 N13508 10
D13508 N13508 0 diode
R13509 N13508 N13509 10
D13509 N13509 0 diode
R13510 N13509 N13510 10
D13510 N13510 0 diode
R13511 N13510 N13511 10
D13511 N13511 0 diode
R13512 N13511 N13512 10
D13512 N13512 0 diode
R13513 N13512 N13513 10
D13513 N13513 0 diode
R13514 N13513 N13514 10
D13514 N13514 0 diode
R13515 N13514 N13515 10
D13515 N13515 0 diode
R13516 N13515 N13516 10
D13516 N13516 0 diode
R13517 N13516 N13517 10
D13517 N13517 0 diode
R13518 N13517 N13518 10
D13518 N13518 0 diode
R13519 N13518 N13519 10
D13519 N13519 0 diode
R13520 N13519 N13520 10
D13520 N13520 0 diode
R13521 N13520 N13521 10
D13521 N13521 0 diode
R13522 N13521 N13522 10
D13522 N13522 0 diode
R13523 N13522 N13523 10
D13523 N13523 0 diode
R13524 N13523 N13524 10
D13524 N13524 0 diode
R13525 N13524 N13525 10
D13525 N13525 0 diode
R13526 N13525 N13526 10
D13526 N13526 0 diode
R13527 N13526 N13527 10
D13527 N13527 0 diode
R13528 N13527 N13528 10
D13528 N13528 0 diode
R13529 N13528 N13529 10
D13529 N13529 0 diode
R13530 N13529 N13530 10
D13530 N13530 0 diode
R13531 N13530 N13531 10
D13531 N13531 0 diode
R13532 N13531 N13532 10
D13532 N13532 0 diode
R13533 N13532 N13533 10
D13533 N13533 0 diode
R13534 N13533 N13534 10
D13534 N13534 0 diode
R13535 N13534 N13535 10
D13535 N13535 0 diode
R13536 N13535 N13536 10
D13536 N13536 0 diode
R13537 N13536 N13537 10
D13537 N13537 0 diode
R13538 N13537 N13538 10
D13538 N13538 0 diode
R13539 N13538 N13539 10
D13539 N13539 0 diode
R13540 N13539 N13540 10
D13540 N13540 0 diode
R13541 N13540 N13541 10
D13541 N13541 0 diode
R13542 N13541 N13542 10
D13542 N13542 0 diode
R13543 N13542 N13543 10
D13543 N13543 0 diode
R13544 N13543 N13544 10
D13544 N13544 0 diode
R13545 N13544 N13545 10
D13545 N13545 0 diode
R13546 N13545 N13546 10
D13546 N13546 0 diode
R13547 N13546 N13547 10
D13547 N13547 0 diode
R13548 N13547 N13548 10
D13548 N13548 0 diode
R13549 N13548 N13549 10
D13549 N13549 0 diode
R13550 N13549 N13550 10
D13550 N13550 0 diode
R13551 N13550 N13551 10
D13551 N13551 0 diode
R13552 N13551 N13552 10
D13552 N13552 0 diode
R13553 N13552 N13553 10
D13553 N13553 0 diode
R13554 N13553 N13554 10
D13554 N13554 0 diode
R13555 N13554 N13555 10
D13555 N13555 0 diode
R13556 N13555 N13556 10
D13556 N13556 0 diode
R13557 N13556 N13557 10
D13557 N13557 0 diode
R13558 N13557 N13558 10
D13558 N13558 0 diode
R13559 N13558 N13559 10
D13559 N13559 0 diode
R13560 N13559 N13560 10
D13560 N13560 0 diode
R13561 N13560 N13561 10
D13561 N13561 0 diode
R13562 N13561 N13562 10
D13562 N13562 0 diode
R13563 N13562 N13563 10
D13563 N13563 0 diode
R13564 N13563 N13564 10
D13564 N13564 0 diode
R13565 N13564 N13565 10
D13565 N13565 0 diode
R13566 N13565 N13566 10
D13566 N13566 0 diode
R13567 N13566 N13567 10
D13567 N13567 0 diode
R13568 N13567 N13568 10
D13568 N13568 0 diode
R13569 N13568 N13569 10
D13569 N13569 0 diode
R13570 N13569 N13570 10
D13570 N13570 0 diode
R13571 N13570 N13571 10
D13571 N13571 0 diode
R13572 N13571 N13572 10
D13572 N13572 0 diode
R13573 N13572 N13573 10
D13573 N13573 0 diode
R13574 N13573 N13574 10
D13574 N13574 0 diode
R13575 N13574 N13575 10
D13575 N13575 0 diode
R13576 N13575 N13576 10
D13576 N13576 0 diode
R13577 N13576 N13577 10
D13577 N13577 0 diode
R13578 N13577 N13578 10
D13578 N13578 0 diode
R13579 N13578 N13579 10
D13579 N13579 0 diode
R13580 N13579 N13580 10
D13580 N13580 0 diode
R13581 N13580 N13581 10
D13581 N13581 0 diode
R13582 N13581 N13582 10
D13582 N13582 0 diode
R13583 N13582 N13583 10
D13583 N13583 0 diode
R13584 N13583 N13584 10
D13584 N13584 0 diode
R13585 N13584 N13585 10
D13585 N13585 0 diode
R13586 N13585 N13586 10
D13586 N13586 0 diode
R13587 N13586 N13587 10
D13587 N13587 0 diode
R13588 N13587 N13588 10
D13588 N13588 0 diode
R13589 N13588 N13589 10
D13589 N13589 0 diode
R13590 N13589 N13590 10
D13590 N13590 0 diode
R13591 N13590 N13591 10
D13591 N13591 0 diode
R13592 N13591 N13592 10
D13592 N13592 0 diode
R13593 N13592 N13593 10
D13593 N13593 0 diode
R13594 N13593 N13594 10
D13594 N13594 0 diode
R13595 N13594 N13595 10
D13595 N13595 0 diode
R13596 N13595 N13596 10
D13596 N13596 0 diode
R13597 N13596 N13597 10
D13597 N13597 0 diode
R13598 N13597 N13598 10
D13598 N13598 0 diode
R13599 N13598 N13599 10
D13599 N13599 0 diode
R13600 N13599 N13600 10
D13600 N13600 0 diode
R13601 N13600 N13601 10
D13601 N13601 0 diode
R13602 N13601 N13602 10
D13602 N13602 0 diode
R13603 N13602 N13603 10
D13603 N13603 0 diode
R13604 N13603 N13604 10
D13604 N13604 0 diode
R13605 N13604 N13605 10
D13605 N13605 0 diode
R13606 N13605 N13606 10
D13606 N13606 0 diode
R13607 N13606 N13607 10
D13607 N13607 0 diode
R13608 N13607 N13608 10
D13608 N13608 0 diode
R13609 N13608 N13609 10
D13609 N13609 0 diode
R13610 N13609 N13610 10
D13610 N13610 0 diode
R13611 N13610 N13611 10
D13611 N13611 0 diode
R13612 N13611 N13612 10
D13612 N13612 0 diode
R13613 N13612 N13613 10
D13613 N13613 0 diode
R13614 N13613 N13614 10
D13614 N13614 0 diode
R13615 N13614 N13615 10
D13615 N13615 0 diode
R13616 N13615 N13616 10
D13616 N13616 0 diode
R13617 N13616 N13617 10
D13617 N13617 0 diode
R13618 N13617 N13618 10
D13618 N13618 0 diode
R13619 N13618 N13619 10
D13619 N13619 0 diode
R13620 N13619 N13620 10
D13620 N13620 0 diode
R13621 N13620 N13621 10
D13621 N13621 0 diode
R13622 N13621 N13622 10
D13622 N13622 0 diode
R13623 N13622 N13623 10
D13623 N13623 0 diode
R13624 N13623 N13624 10
D13624 N13624 0 diode
R13625 N13624 N13625 10
D13625 N13625 0 diode
R13626 N13625 N13626 10
D13626 N13626 0 diode
R13627 N13626 N13627 10
D13627 N13627 0 diode
R13628 N13627 N13628 10
D13628 N13628 0 diode
R13629 N13628 N13629 10
D13629 N13629 0 diode
R13630 N13629 N13630 10
D13630 N13630 0 diode
R13631 N13630 N13631 10
D13631 N13631 0 diode
R13632 N13631 N13632 10
D13632 N13632 0 diode
R13633 N13632 N13633 10
D13633 N13633 0 diode
R13634 N13633 N13634 10
D13634 N13634 0 diode
R13635 N13634 N13635 10
D13635 N13635 0 diode
R13636 N13635 N13636 10
D13636 N13636 0 diode
R13637 N13636 N13637 10
D13637 N13637 0 diode
R13638 N13637 N13638 10
D13638 N13638 0 diode
R13639 N13638 N13639 10
D13639 N13639 0 diode
R13640 N13639 N13640 10
D13640 N13640 0 diode
R13641 N13640 N13641 10
D13641 N13641 0 diode
R13642 N13641 N13642 10
D13642 N13642 0 diode
R13643 N13642 N13643 10
D13643 N13643 0 diode
R13644 N13643 N13644 10
D13644 N13644 0 diode
R13645 N13644 N13645 10
D13645 N13645 0 diode
R13646 N13645 N13646 10
D13646 N13646 0 diode
R13647 N13646 N13647 10
D13647 N13647 0 diode
R13648 N13647 N13648 10
D13648 N13648 0 diode
R13649 N13648 N13649 10
D13649 N13649 0 diode
R13650 N13649 N13650 10
D13650 N13650 0 diode
R13651 N13650 N13651 10
D13651 N13651 0 diode
R13652 N13651 N13652 10
D13652 N13652 0 diode
R13653 N13652 N13653 10
D13653 N13653 0 diode
R13654 N13653 N13654 10
D13654 N13654 0 diode
R13655 N13654 N13655 10
D13655 N13655 0 diode
R13656 N13655 N13656 10
D13656 N13656 0 diode
R13657 N13656 N13657 10
D13657 N13657 0 diode
R13658 N13657 N13658 10
D13658 N13658 0 diode
R13659 N13658 N13659 10
D13659 N13659 0 diode
R13660 N13659 N13660 10
D13660 N13660 0 diode
R13661 N13660 N13661 10
D13661 N13661 0 diode
R13662 N13661 N13662 10
D13662 N13662 0 diode
R13663 N13662 N13663 10
D13663 N13663 0 diode
R13664 N13663 N13664 10
D13664 N13664 0 diode
R13665 N13664 N13665 10
D13665 N13665 0 diode
R13666 N13665 N13666 10
D13666 N13666 0 diode
R13667 N13666 N13667 10
D13667 N13667 0 diode
R13668 N13667 N13668 10
D13668 N13668 0 diode
R13669 N13668 N13669 10
D13669 N13669 0 diode
R13670 N13669 N13670 10
D13670 N13670 0 diode
R13671 N13670 N13671 10
D13671 N13671 0 diode
R13672 N13671 N13672 10
D13672 N13672 0 diode
R13673 N13672 N13673 10
D13673 N13673 0 diode
R13674 N13673 N13674 10
D13674 N13674 0 diode
R13675 N13674 N13675 10
D13675 N13675 0 diode
R13676 N13675 N13676 10
D13676 N13676 0 diode
R13677 N13676 N13677 10
D13677 N13677 0 diode
R13678 N13677 N13678 10
D13678 N13678 0 diode
R13679 N13678 N13679 10
D13679 N13679 0 diode
R13680 N13679 N13680 10
D13680 N13680 0 diode
R13681 N13680 N13681 10
D13681 N13681 0 diode
R13682 N13681 N13682 10
D13682 N13682 0 diode
R13683 N13682 N13683 10
D13683 N13683 0 diode
R13684 N13683 N13684 10
D13684 N13684 0 diode
R13685 N13684 N13685 10
D13685 N13685 0 diode
R13686 N13685 N13686 10
D13686 N13686 0 diode
R13687 N13686 N13687 10
D13687 N13687 0 diode
R13688 N13687 N13688 10
D13688 N13688 0 diode
R13689 N13688 N13689 10
D13689 N13689 0 diode
R13690 N13689 N13690 10
D13690 N13690 0 diode
R13691 N13690 N13691 10
D13691 N13691 0 diode
R13692 N13691 N13692 10
D13692 N13692 0 diode
R13693 N13692 N13693 10
D13693 N13693 0 diode
R13694 N13693 N13694 10
D13694 N13694 0 diode
R13695 N13694 N13695 10
D13695 N13695 0 diode
R13696 N13695 N13696 10
D13696 N13696 0 diode
R13697 N13696 N13697 10
D13697 N13697 0 diode
R13698 N13697 N13698 10
D13698 N13698 0 diode
R13699 N13698 N13699 10
D13699 N13699 0 diode
R13700 N13699 N13700 10
D13700 N13700 0 diode
R13701 N13700 N13701 10
D13701 N13701 0 diode
R13702 N13701 N13702 10
D13702 N13702 0 diode
R13703 N13702 N13703 10
D13703 N13703 0 diode
R13704 N13703 N13704 10
D13704 N13704 0 diode
R13705 N13704 N13705 10
D13705 N13705 0 diode
R13706 N13705 N13706 10
D13706 N13706 0 diode
R13707 N13706 N13707 10
D13707 N13707 0 diode
R13708 N13707 N13708 10
D13708 N13708 0 diode
R13709 N13708 N13709 10
D13709 N13709 0 diode
R13710 N13709 N13710 10
D13710 N13710 0 diode
R13711 N13710 N13711 10
D13711 N13711 0 diode
R13712 N13711 N13712 10
D13712 N13712 0 diode
R13713 N13712 N13713 10
D13713 N13713 0 diode
R13714 N13713 N13714 10
D13714 N13714 0 diode
R13715 N13714 N13715 10
D13715 N13715 0 diode
R13716 N13715 N13716 10
D13716 N13716 0 diode
R13717 N13716 N13717 10
D13717 N13717 0 diode
R13718 N13717 N13718 10
D13718 N13718 0 diode
R13719 N13718 N13719 10
D13719 N13719 0 diode
R13720 N13719 N13720 10
D13720 N13720 0 diode
R13721 N13720 N13721 10
D13721 N13721 0 diode
R13722 N13721 N13722 10
D13722 N13722 0 diode
R13723 N13722 N13723 10
D13723 N13723 0 diode
R13724 N13723 N13724 10
D13724 N13724 0 diode
R13725 N13724 N13725 10
D13725 N13725 0 diode
R13726 N13725 N13726 10
D13726 N13726 0 diode
R13727 N13726 N13727 10
D13727 N13727 0 diode
R13728 N13727 N13728 10
D13728 N13728 0 diode
R13729 N13728 N13729 10
D13729 N13729 0 diode
R13730 N13729 N13730 10
D13730 N13730 0 diode
R13731 N13730 N13731 10
D13731 N13731 0 diode
R13732 N13731 N13732 10
D13732 N13732 0 diode
R13733 N13732 N13733 10
D13733 N13733 0 diode
R13734 N13733 N13734 10
D13734 N13734 0 diode
R13735 N13734 N13735 10
D13735 N13735 0 diode
R13736 N13735 N13736 10
D13736 N13736 0 diode
R13737 N13736 N13737 10
D13737 N13737 0 diode
R13738 N13737 N13738 10
D13738 N13738 0 diode
R13739 N13738 N13739 10
D13739 N13739 0 diode
R13740 N13739 N13740 10
D13740 N13740 0 diode
R13741 N13740 N13741 10
D13741 N13741 0 diode
R13742 N13741 N13742 10
D13742 N13742 0 diode
R13743 N13742 N13743 10
D13743 N13743 0 diode
R13744 N13743 N13744 10
D13744 N13744 0 diode
R13745 N13744 N13745 10
D13745 N13745 0 diode
R13746 N13745 N13746 10
D13746 N13746 0 diode
R13747 N13746 N13747 10
D13747 N13747 0 diode
R13748 N13747 N13748 10
D13748 N13748 0 diode
R13749 N13748 N13749 10
D13749 N13749 0 diode
R13750 N13749 N13750 10
D13750 N13750 0 diode
R13751 N13750 N13751 10
D13751 N13751 0 diode
R13752 N13751 N13752 10
D13752 N13752 0 diode
R13753 N13752 N13753 10
D13753 N13753 0 diode
R13754 N13753 N13754 10
D13754 N13754 0 diode
R13755 N13754 N13755 10
D13755 N13755 0 diode
R13756 N13755 N13756 10
D13756 N13756 0 diode
R13757 N13756 N13757 10
D13757 N13757 0 diode
R13758 N13757 N13758 10
D13758 N13758 0 diode
R13759 N13758 N13759 10
D13759 N13759 0 diode
R13760 N13759 N13760 10
D13760 N13760 0 diode
R13761 N13760 N13761 10
D13761 N13761 0 diode
R13762 N13761 N13762 10
D13762 N13762 0 diode
R13763 N13762 N13763 10
D13763 N13763 0 diode
R13764 N13763 N13764 10
D13764 N13764 0 diode
R13765 N13764 N13765 10
D13765 N13765 0 diode
R13766 N13765 N13766 10
D13766 N13766 0 diode
R13767 N13766 N13767 10
D13767 N13767 0 diode
R13768 N13767 N13768 10
D13768 N13768 0 diode
R13769 N13768 N13769 10
D13769 N13769 0 diode
R13770 N13769 N13770 10
D13770 N13770 0 diode
R13771 N13770 N13771 10
D13771 N13771 0 diode
R13772 N13771 N13772 10
D13772 N13772 0 diode
R13773 N13772 N13773 10
D13773 N13773 0 diode
R13774 N13773 N13774 10
D13774 N13774 0 diode
R13775 N13774 N13775 10
D13775 N13775 0 diode
R13776 N13775 N13776 10
D13776 N13776 0 diode
R13777 N13776 N13777 10
D13777 N13777 0 diode
R13778 N13777 N13778 10
D13778 N13778 0 diode
R13779 N13778 N13779 10
D13779 N13779 0 diode
R13780 N13779 N13780 10
D13780 N13780 0 diode
R13781 N13780 N13781 10
D13781 N13781 0 diode
R13782 N13781 N13782 10
D13782 N13782 0 diode
R13783 N13782 N13783 10
D13783 N13783 0 diode
R13784 N13783 N13784 10
D13784 N13784 0 diode
R13785 N13784 N13785 10
D13785 N13785 0 diode
R13786 N13785 N13786 10
D13786 N13786 0 diode
R13787 N13786 N13787 10
D13787 N13787 0 diode
R13788 N13787 N13788 10
D13788 N13788 0 diode
R13789 N13788 N13789 10
D13789 N13789 0 diode
R13790 N13789 N13790 10
D13790 N13790 0 diode
R13791 N13790 N13791 10
D13791 N13791 0 diode
R13792 N13791 N13792 10
D13792 N13792 0 diode
R13793 N13792 N13793 10
D13793 N13793 0 diode
R13794 N13793 N13794 10
D13794 N13794 0 diode
R13795 N13794 N13795 10
D13795 N13795 0 diode
R13796 N13795 N13796 10
D13796 N13796 0 diode
R13797 N13796 N13797 10
D13797 N13797 0 diode
R13798 N13797 N13798 10
D13798 N13798 0 diode
R13799 N13798 N13799 10
D13799 N13799 0 diode
R13800 N13799 N13800 10
D13800 N13800 0 diode
R13801 N13800 N13801 10
D13801 N13801 0 diode
R13802 N13801 N13802 10
D13802 N13802 0 diode
R13803 N13802 N13803 10
D13803 N13803 0 diode
R13804 N13803 N13804 10
D13804 N13804 0 diode
R13805 N13804 N13805 10
D13805 N13805 0 diode
R13806 N13805 N13806 10
D13806 N13806 0 diode
R13807 N13806 N13807 10
D13807 N13807 0 diode
R13808 N13807 N13808 10
D13808 N13808 0 diode
R13809 N13808 N13809 10
D13809 N13809 0 diode
R13810 N13809 N13810 10
D13810 N13810 0 diode
R13811 N13810 N13811 10
D13811 N13811 0 diode
R13812 N13811 N13812 10
D13812 N13812 0 diode
R13813 N13812 N13813 10
D13813 N13813 0 diode
R13814 N13813 N13814 10
D13814 N13814 0 diode
R13815 N13814 N13815 10
D13815 N13815 0 diode
R13816 N13815 N13816 10
D13816 N13816 0 diode
R13817 N13816 N13817 10
D13817 N13817 0 diode
R13818 N13817 N13818 10
D13818 N13818 0 diode
R13819 N13818 N13819 10
D13819 N13819 0 diode
R13820 N13819 N13820 10
D13820 N13820 0 diode
R13821 N13820 N13821 10
D13821 N13821 0 diode
R13822 N13821 N13822 10
D13822 N13822 0 diode
R13823 N13822 N13823 10
D13823 N13823 0 diode
R13824 N13823 N13824 10
D13824 N13824 0 diode
R13825 N13824 N13825 10
D13825 N13825 0 diode
R13826 N13825 N13826 10
D13826 N13826 0 diode
R13827 N13826 N13827 10
D13827 N13827 0 diode
R13828 N13827 N13828 10
D13828 N13828 0 diode
R13829 N13828 N13829 10
D13829 N13829 0 diode
R13830 N13829 N13830 10
D13830 N13830 0 diode
R13831 N13830 N13831 10
D13831 N13831 0 diode
R13832 N13831 N13832 10
D13832 N13832 0 diode
R13833 N13832 N13833 10
D13833 N13833 0 diode
R13834 N13833 N13834 10
D13834 N13834 0 diode
R13835 N13834 N13835 10
D13835 N13835 0 diode
R13836 N13835 N13836 10
D13836 N13836 0 diode
R13837 N13836 N13837 10
D13837 N13837 0 diode
R13838 N13837 N13838 10
D13838 N13838 0 diode
R13839 N13838 N13839 10
D13839 N13839 0 diode
R13840 N13839 N13840 10
D13840 N13840 0 diode
R13841 N13840 N13841 10
D13841 N13841 0 diode
R13842 N13841 N13842 10
D13842 N13842 0 diode
R13843 N13842 N13843 10
D13843 N13843 0 diode
R13844 N13843 N13844 10
D13844 N13844 0 diode
R13845 N13844 N13845 10
D13845 N13845 0 diode
R13846 N13845 N13846 10
D13846 N13846 0 diode
R13847 N13846 N13847 10
D13847 N13847 0 diode
R13848 N13847 N13848 10
D13848 N13848 0 diode
R13849 N13848 N13849 10
D13849 N13849 0 diode
R13850 N13849 N13850 10
D13850 N13850 0 diode
R13851 N13850 N13851 10
D13851 N13851 0 diode
R13852 N13851 N13852 10
D13852 N13852 0 diode
R13853 N13852 N13853 10
D13853 N13853 0 diode
R13854 N13853 N13854 10
D13854 N13854 0 diode
R13855 N13854 N13855 10
D13855 N13855 0 diode
R13856 N13855 N13856 10
D13856 N13856 0 diode
R13857 N13856 N13857 10
D13857 N13857 0 diode
R13858 N13857 N13858 10
D13858 N13858 0 diode
R13859 N13858 N13859 10
D13859 N13859 0 diode
R13860 N13859 N13860 10
D13860 N13860 0 diode
R13861 N13860 N13861 10
D13861 N13861 0 diode
R13862 N13861 N13862 10
D13862 N13862 0 diode
R13863 N13862 N13863 10
D13863 N13863 0 diode
R13864 N13863 N13864 10
D13864 N13864 0 diode
R13865 N13864 N13865 10
D13865 N13865 0 diode
R13866 N13865 N13866 10
D13866 N13866 0 diode
R13867 N13866 N13867 10
D13867 N13867 0 diode
R13868 N13867 N13868 10
D13868 N13868 0 diode
R13869 N13868 N13869 10
D13869 N13869 0 diode
R13870 N13869 N13870 10
D13870 N13870 0 diode
R13871 N13870 N13871 10
D13871 N13871 0 diode
R13872 N13871 N13872 10
D13872 N13872 0 diode
R13873 N13872 N13873 10
D13873 N13873 0 diode
R13874 N13873 N13874 10
D13874 N13874 0 diode
R13875 N13874 N13875 10
D13875 N13875 0 diode
R13876 N13875 N13876 10
D13876 N13876 0 diode
R13877 N13876 N13877 10
D13877 N13877 0 diode
R13878 N13877 N13878 10
D13878 N13878 0 diode
R13879 N13878 N13879 10
D13879 N13879 0 diode
R13880 N13879 N13880 10
D13880 N13880 0 diode
R13881 N13880 N13881 10
D13881 N13881 0 diode
R13882 N13881 N13882 10
D13882 N13882 0 diode
R13883 N13882 N13883 10
D13883 N13883 0 diode
R13884 N13883 N13884 10
D13884 N13884 0 diode
R13885 N13884 N13885 10
D13885 N13885 0 diode
R13886 N13885 N13886 10
D13886 N13886 0 diode
R13887 N13886 N13887 10
D13887 N13887 0 diode
R13888 N13887 N13888 10
D13888 N13888 0 diode
R13889 N13888 N13889 10
D13889 N13889 0 diode
R13890 N13889 N13890 10
D13890 N13890 0 diode
R13891 N13890 N13891 10
D13891 N13891 0 diode
R13892 N13891 N13892 10
D13892 N13892 0 diode
R13893 N13892 N13893 10
D13893 N13893 0 diode
R13894 N13893 N13894 10
D13894 N13894 0 diode
R13895 N13894 N13895 10
D13895 N13895 0 diode
R13896 N13895 N13896 10
D13896 N13896 0 diode
R13897 N13896 N13897 10
D13897 N13897 0 diode
R13898 N13897 N13898 10
D13898 N13898 0 diode
R13899 N13898 N13899 10
D13899 N13899 0 diode
R13900 N13899 N13900 10
D13900 N13900 0 diode
R13901 N13900 N13901 10
D13901 N13901 0 diode
R13902 N13901 N13902 10
D13902 N13902 0 diode
R13903 N13902 N13903 10
D13903 N13903 0 diode
R13904 N13903 N13904 10
D13904 N13904 0 diode
R13905 N13904 N13905 10
D13905 N13905 0 diode
R13906 N13905 N13906 10
D13906 N13906 0 diode
R13907 N13906 N13907 10
D13907 N13907 0 diode
R13908 N13907 N13908 10
D13908 N13908 0 diode
R13909 N13908 N13909 10
D13909 N13909 0 diode
R13910 N13909 N13910 10
D13910 N13910 0 diode
R13911 N13910 N13911 10
D13911 N13911 0 diode
R13912 N13911 N13912 10
D13912 N13912 0 diode
R13913 N13912 N13913 10
D13913 N13913 0 diode
R13914 N13913 N13914 10
D13914 N13914 0 diode
R13915 N13914 N13915 10
D13915 N13915 0 diode
R13916 N13915 N13916 10
D13916 N13916 0 diode
R13917 N13916 N13917 10
D13917 N13917 0 diode
R13918 N13917 N13918 10
D13918 N13918 0 diode
R13919 N13918 N13919 10
D13919 N13919 0 diode
R13920 N13919 N13920 10
D13920 N13920 0 diode
R13921 N13920 N13921 10
D13921 N13921 0 diode
R13922 N13921 N13922 10
D13922 N13922 0 diode
R13923 N13922 N13923 10
D13923 N13923 0 diode
R13924 N13923 N13924 10
D13924 N13924 0 diode
R13925 N13924 N13925 10
D13925 N13925 0 diode
R13926 N13925 N13926 10
D13926 N13926 0 diode
R13927 N13926 N13927 10
D13927 N13927 0 diode
R13928 N13927 N13928 10
D13928 N13928 0 diode
R13929 N13928 N13929 10
D13929 N13929 0 diode
R13930 N13929 N13930 10
D13930 N13930 0 diode
R13931 N13930 N13931 10
D13931 N13931 0 diode
R13932 N13931 N13932 10
D13932 N13932 0 diode
R13933 N13932 N13933 10
D13933 N13933 0 diode
R13934 N13933 N13934 10
D13934 N13934 0 diode
R13935 N13934 N13935 10
D13935 N13935 0 diode
R13936 N13935 N13936 10
D13936 N13936 0 diode
R13937 N13936 N13937 10
D13937 N13937 0 diode
R13938 N13937 N13938 10
D13938 N13938 0 diode
R13939 N13938 N13939 10
D13939 N13939 0 diode
R13940 N13939 N13940 10
D13940 N13940 0 diode
R13941 N13940 N13941 10
D13941 N13941 0 diode
R13942 N13941 N13942 10
D13942 N13942 0 diode
R13943 N13942 N13943 10
D13943 N13943 0 diode
R13944 N13943 N13944 10
D13944 N13944 0 diode
R13945 N13944 N13945 10
D13945 N13945 0 diode
R13946 N13945 N13946 10
D13946 N13946 0 diode
R13947 N13946 N13947 10
D13947 N13947 0 diode
R13948 N13947 N13948 10
D13948 N13948 0 diode
R13949 N13948 N13949 10
D13949 N13949 0 diode
R13950 N13949 N13950 10
D13950 N13950 0 diode
R13951 N13950 N13951 10
D13951 N13951 0 diode
R13952 N13951 N13952 10
D13952 N13952 0 diode
R13953 N13952 N13953 10
D13953 N13953 0 diode
R13954 N13953 N13954 10
D13954 N13954 0 diode
R13955 N13954 N13955 10
D13955 N13955 0 diode
R13956 N13955 N13956 10
D13956 N13956 0 diode
R13957 N13956 N13957 10
D13957 N13957 0 diode
R13958 N13957 N13958 10
D13958 N13958 0 diode
R13959 N13958 N13959 10
D13959 N13959 0 diode
R13960 N13959 N13960 10
D13960 N13960 0 diode
R13961 N13960 N13961 10
D13961 N13961 0 diode
R13962 N13961 N13962 10
D13962 N13962 0 diode
R13963 N13962 N13963 10
D13963 N13963 0 diode
R13964 N13963 N13964 10
D13964 N13964 0 diode
R13965 N13964 N13965 10
D13965 N13965 0 diode
R13966 N13965 N13966 10
D13966 N13966 0 diode
R13967 N13966 N13967 10
D13967 N13967 0 diode
R13968 N13967 N13968 10
D13968 N13968 0 diode
R13969 N13968 N13969 10
D13969 N13969 0 diode
R13970 N13969 N13970 10
D13970 N13970 0 diode
R13971 N13970 N13971 10
D13971 N13971 0 diode
R13972 N13971 N13972 10
D13972 N13972 0 diode
R13973 N13972 N13973 10
D13973 N13973 0 diode
R13974 N13973 N13974 10
D13974 N13974 0 diode
R13975 N13974 N13975 10
D13975 N13975 0 diode
R13976 N13975 N13976 10
D13976 N13976 0 diode
R13977 N13976 N13977 10
D13977 N13977 0 diode
R13978 N13977 N13978 10
D13978 N13978 0 diode
R13979 N13978 N13979 10
D13979 N13979 0 diode
R13980 N13979 N13980 10
D13980 N13980 0 diode
R13981 N13980 N13981 10
D13981 N13981 0 diode
R13982 N13981 N13982 10
D13982 N13982 0 diode
R13983 N13982 N13983 10
D13983 N13983 0 diode
R13984 N13983 N13984 10
D13984 N13984 0 diode
R13985 N13984 N13985 10
D13985 N13985 0 diode
R13986 N13985 N13986 10
D13986 N13986 0 diode
R13987 N13986 N13987 10
D13987 N13987 0 diode
R13988 N13987 N13988 10
D13988 N13988 0 diode
R13989 N13988 N13989 10
D13989 N13989 0 diode
R13990 N13989 N13990 10
D13990 N13990 0 diode
R13991 N13990 N13991 10
D13991 N13991 0 diode
R13992 N13991 N13992 10
D13992 N13992 0 diode
R13993 N13992 N13993 10
D13993 N13993 0 diode
R13994 N13993 N13994 10
D13994 N13994 0 diode
R13995 N13994 N13995 10
D13995 N13995 0 diode
R13996 N13995 N13996 10
D13996 N13996 0 diode
R13997 N13996 N13997 10
D13997 N13997 0 diode
R13998 N13997 N13998 10
D13998 N13998 0 diode
R13999 N13998 N13999 10
D13999 N13999 0 diode
R14000 N13999 N14000 10
D14000 N14000 0 diode
R14001 N14000 N14001 10
D14001 N14001 0 diode
R14002 N14001 N14002 10
D14002 N14002 0 diode
R14003 N14002 N14003 10
D14003 N14003 0 diode
R14004 N14003 N14004 10
D14004 N14004 0 diode
R14005 N14004 N14005 10
D14005 N14005 0 diode
R14006 N14005 N14006 10
D14006 N14006 0 diode
R14007 N14006 N14007 10
D14007 N14007 0 diode
R14008 N14007 N14008 10
D14008 N14008 0 diode
R14009 N14008 N14009 10
D14009 N14009 0 diode
R14010 N14009 N14010 10
D14010 N14010 0 diode
R14011 N14010 N14011 10
D14011 N14011 0 diode
R14012 N14011 N14012 10
D14012 N14012 0 diode
R14013 N14012 N14013 10
D14013 N14013 0 diode
R14014 N14013 N14014 10
D14014 N14014 0 diode
R14015 N14014 N14015 10
D14015 N14015 0 diode
R14016 N14015 N14016 10
D14016 N14016 0 diode
R14017 N14016 N14017 10
D14017 N14017 0 diode
R14018 N14017 N14018 10
D14018 N14018 0 diode
R14019 N14018 N14019 10
D14019 N14019 0 diode
R14020 N14019 N14020 10
D14020 N14020 0 diode
R14021 N14020 N14021 10
D14021 N14021 0 diode
R14022 N14021 N14022 10
D14022 N14022 0 diode
R14023 N14022 N14023 10
D14023 N14023 0 diode
R14024 N14023 N14024 10
D14024 N14024 0 diode
R14025 N14024 N14025 10
D14025 N14025 0 diode
R14026 N14025 N14026 10
D14026 N14026 0 diode
R14027 N14026 N14027 10
D14027 N14027 0 diode
R14028 N14027 N14028 10
D14028 N14028 0 diode
R14029 N14028 N14029 10
D14029 N14029 0 diode
R14030 N14029 N14030 10
D14030 N14030 0 diode
R14031 N14030 N14031 10
D14031 N14031 0 diode
R14032 N14031 N14032 10
D14032 N14032 0 diode
R14033 N14032 N14033 10
D14033 N14033 0 diode
R14034 N14033 N14034 10
D14034 N14034 0 diode
R14035 N14034 N14035 10
D14035 N14035 0 diode
R14036 N14035 N14036 10
D14036 N14036 0 diode
R14037 N14036 N14037 10
D14037 N14037 0 diode
R14038 N14037 N14038 10
D14038 N14038 0 diode
R14039 N14038 N14039 10
D14039 N14039 0 diode
R14040 N14039 N14040 10
D14040 N14040 0 diode
R14041 N14040 N14041 10
D14041 N14041 0 diode
R14042 N14041 N14042 10
D14042 N14042 0 diode
R14043 N14042 N14043 10
D14043 N14043 0 diode
R14044 N14043 N14044 10
D14044 N14044 0 diode
R14045 N14044 N14045 10
D14045 N14045 0 diode
R14046 N14045 N14046 10
D14046 N14046 0 diode
R14047 N14046 N14047 10
D14047 N14047 0 diode
R14048 N14047 N14048 10
D14048 N14048 0 diode
R14049 N14048 N14049 10
D14049 N14049 0 diode
R14050 N14049 N14050 10
D14050 N14050 0 diode
R14051 N14050 N14051 10
D14051 N14051 0 diode
R14052 N14051 N14052 10
D14052 N14052 0 diode
R14053 N14052 N14053 10
D14053 N14053 0 diode
R14054 N14053 N14054 10
D14054 N14054 0 diode
R14055 N14054 N14055 10
D14055 N14055 0 diode
R14056 N14055 N14056 10
D14056 N14056 0 diode
R14057 N14056 N14057 10
D14057 N14057 0 diode
R14058 N14057 N14058 10
D14058 N14058 0 diode
R14059 N14058 N14059 10
D14059 N14059 0 diode
R14060 N14059 N14060 10
D14060 N14060 0 diode
R14061 N14060 N14061 10
D14061 N14061 0 diode
R14062 N14061 N14062 10
D14062 N14062 0 diode
R14063 N14062 N14063 10
D14063 N14063 0 diode
R14064 N14063 N14064 10
D14064 N14064 0 diode
R14065 N14064 N14065 10
D14065 N14065 0 diode
R14066 N14065 N14066 10
D14066 N14066 0 diode
R14067 N14066 N14067 10
D14067 N14067 0 diode
R14068 N14067 N14068 10
D14068 N14068 0 diode
R14069 N14068 N14069 10
D14069 N14069 0 diode
R14070 N14069 N14070 10
D14070 N14070 0 diode
R14071 N14070 N14071 10
D14071 N14071 0 diode
R14072 N14071 N14072 10
D14072 N14072 0 diode
R14073 N14072 N14073 10
D14073 N14073 0 diode
R14074 N14073 N14074 10
D14074 N14074 0 diode
R14075 N14074 N14075 10
D14075 N14075 0 diode
R14076 N14075 N14076 10
D14076 N14076 0 diode
R14077 N14076 N14077 10
D14077 N14077 0 diode
R14078 N14077 N14078 10
D14078 N14078 0 diode
R14079 N14078 N14079 10
D14079 N14079 0 diode
R14080 N14079 N14080 10
D14080 N14080 0 diode
R14081 N14080 N14081 10
D14081 N14081 0 diode
R14082 N14081 N14082 10
D14082 N14082 0 diode
R14083 N14082 N14083 10
D14083 N14083 0 diode
R14084 N14083 N14084 10
D14084 N14084 0 diode
R14085 N14084 N14085 10
D14085 N14085 0 diode
R14086 N14085 N14086 10
D14086 N14086 0 diode
R14087 N14086 N14087 10
D14087 N14087 0 diode
R14088 N14087 N14088 10
D14088 N14088 0 diode
R14089 N14088 N14089 10
D14089 N14089 0 diode
R14090 N14089 N14090 10
D14090 N14090 0 diode
R14091 N14090 N14091 10
D14091 N14091 0 diode
R14092 N14091 N14092 10
D14092 N14092 0 diode
R14093 N14092 N14093 10
D14093 N14093 0 diode
R14094 N14093 N14094 10
D14094 N14094 0 diode
R14095 N14094 N14095 10
D14095 N14095 0 diode
R14096 N14095 N14096 10
D14096 N14096 0 diode
R14097 N14096 N14097 10
D14097 N14097 0 diode
R14098 N14097 N14098 10
D14098 N14098 0 diode
R14099 N14098 N14099 10
D14099 N14099 0 diode
R14100 N14099 N14100 10
D14100 N14100 0 diode
R14101 N14100 N14101 10
D14101 N14101 0 diode
R14102 N14101 N14102 10
D14102 N14102 0 diode
R14103 N14102 N14103 10
D14103 N14103 0 diode
R14104 N14103 N14104 10
D14104 N14104 0 diode
R14105 N14104 N14105 10
D14105 N14105 0 diode
R14106 N14105 N14106 10
D14106 N14106 0 diode
R14107 N14106 N14107 10
D14107 N14107 0 diode
R14108 N14107 N14108 10
D14108 N14108 0 diode
R14109 N14108 N14109 10
D14109 N14109 0 diode
R14110 N14109 N14110 10
D14110 N14110 0 diode
R14111 N14110 N14111 10
D14111 N14111 0 diode
R14112 N14111 N14112 10
D14112 N14112 0 diode
R14113 N14112 N14113 10
D14113 N14113 0 diode
R14114 N14113 N14114 10
D14114 N14114 0 diode
R14115 N14114 N14115 10
D14115 N14115 0 diode
R14116 N14115 N14116 10
D14116 N14116 0 diode
R14117 N14116 N14117 10
D14117 N14117 0 diode
R14118 N14117 N14118 10
D14118 N14118 0 diode
R14119 N14118 N14119 10
D14119 N14119 0 diode
R14120 N14119 N14120 10
D14120 N14120 0 diode
R14121 N14120 N14121 10
D14121 N14121 0 diode
R14122 N14121 N14122 10
D14122 N14122 0 diode
R14123 N14122 N14123 10
D14123 N14123 0 diode
R14124 N14123 N14124 10
D14124 N14124 0 diode
R14125 N14124 N14125 10
D14125 N14125 0 diode
R14126 N14125 N14126 10
D14126 N14126 0 diode
R14127 N14126 N14127 10
D14127 N14127 0 diode
R14128 N14127 N14128 10
D14128 N14128 0 diode
R14129 N14128 N14129 10
D14129 N14129 0 diode
R14130 N14129 N14130 10
D14130 N14130 0 diode
R14131 N14130 N14131 10
D14131 N14131 0 diode
R14132 N14131 N14132 10
D14132 N14132 0 diode
R14133 N14132 N14133 10
D14133 N14133 0 diode
R14134 N14133 N14134 10
D14134 N14134 0 diode
R14135 N14134 N14135 10
D14135 N14135 0 diode
R14136 N14135 N14136 10
D14136 N14136 0 diode
R14137 N14136 N14137 10
D14137 N14137 0 diode
R14138 N14137 N14138 10
D14138 N14138 0 diode
R14139 N14138 N14139 10
D14139 N14139 0 diode
R14140 N14139 N14140 10
D14140 N14140 0 diode
R14141 N14140 N14141 10
D14141 N14141 0 diode
R14142 N14141 N14142 10
D14142 N14142 0 diode
R14143 N14142 N14143 10
D14143 N14143 0 diode
R14144 N14143 N14144 10
D14144 N14144 0 diode
R14145 N14144 N14145 10
D14145 N14145 0 diode
R14146 N14145 N14146 10
D14146 N14146 0 diode
R14147 N14146 N14147 10
D14147 N14147 0 diode
R14148 N14147 N14148 10
D14148 N14148 0 diode
R14149 N14148 N14149 10
D14149 N14149 0 diode
R14150 N14149 N14150 10
D14150 N14150 0 diode
R14151 N14150 N14151 10
D14151 N14151 0 diode
R14152 N14151 N14152 10
D14152 N14152 0 diode
R14153 N14152 N14153 10
D14153 N14153 0 diode
R14154 N14153 N14154 10
D14154 N14154 0 diode
R14155 N14154 N14155 10
D14155 N14155 0 diode
R14156 N14155 N14156 10
D14156 N14156 0 diode
R14157 N14156 N14157 10
D14157 N14157 0 diode
R14158 N14157 N14158 10
D14158 N14158 0 diode
R14159 N14158 N14159 10
D14159 N14159 0 diode
R14160 N14159 N14160 10
D14160 N14160 0 diode
R14161 N14160 N14161 10
D14161 N14161 0 diode
R14162 N14161 N14162 10
D14162 N14162 0 diode
R14163 N14162 N14163 10
D14163 N14163 0 diode
R14164 N14163 N14164 10
D14164 N14164 0 diode
R14165 N14164 N14165 10
D14165 N14165 0 diode
R14166 N14165 N14166 10
D14166 N14166 0 diode
R14167 N14166 N14167 10
D14167 N14167 0 diode
R14168 N14167 N14168 10
D14168 N14168 0 diode
R14169 N14168 N14169 10
D14169 N14169 0 diode
R14170 N14169 N14170 10
D14170 N14170 0 diode
R14171 N14170 N14171 10
D14171 N14171 0 diode
R14172 N14171 N14172 10
D14172 N14172 0 diode
R14173 N14172 N14173 10
D14173 N14173 0 diode
R14174 N14173 N14174 10
D14174 N14174 0 diode
R14175 N14174 N14175 10
D14175 N14175 0 diode
R14176 N14175 N14176 10
D14176 N14176 0 diode
R14177 N14176 N14177 10
D14177 N14177 0 diode
R14178 N14177 N14178 10
D14178 N14178 0 diode
R14179 N14178 N14179 10
D14179 N14179 0 diode
R14180 N14179 N14180 10
D14180 N14180 0 diode
R14181 N14180 N14181 10
D14181 N14181 0 diode
R14182 N14181 N14182 10
D14182 N14182 0 diode
R14183 N14182 N14183 10
D14183 N14183 0 diode
R14184 N14183 N14184 10
D14184 N14184 0 diode
R14185 N14184 N14185 10
D14185 N14185 0 diode
R14186 N14185 N14186 10
D14186 N14186 0 diode
R14187 N14186 N14187 10
D14187 N14187 0 diode
R14188 N14187 N14188 10
D14188 N14188 0 diode
R14189 N14188 N14189 10
D14189 N14189 0 diode
R14190 N14189 N14190 10
D14190 N14190 0 diode
R14191 N14190 N14191 10
D14191 N14191 0 diode
R14192 N14191 N14192 10
D14192 N14192 0 diode
R14193 N14192 N14193 10
D14193 N14193 0 diode
R14194 N14193 N14194 10
D14194 N14194 0 diode
R14195 N14194 N14195 10
D14195 N14195 0 diode
R14196 N14195 N14196 10
D14196 N14196 0 diode
R14197 N14196 N14197 10
D14197 N14197 0 diode
R14198 N14197 N14198 10
D14198 N14198 0 diode
R14199 N14198 N14199 10
D14199 N14199 0 diode
R14200 N14199 N14200 10
D14200 N14200 0 diode
R14201 N14200 N14201 10
D14201 N14201 0 diode
R14202 N14201 N14202 10
D14202 N14202 0 diode
R14203 N14202 N14203 10
D14203 N14203 0 diode
R14204 N14203 N14204 10
D14204 N14204 0 diode
R14205 N14204 N14205 10
D14205 N14205 0 diode
R14206 N14205 N14206 10
D14206 N14206 0 diode
R14207 N14206 N14207 10
D14207 N14207 0 diode
R14208 N14207 N14208 10
D14208 N14208 0 diode
R14209 N14208 N14209 10
D14209 N14209 0 diode
R14210 N14209 N14210 10
D14210 N14210 0 diode
R14211 N14210 N14211 10
D14211 N14211 0 diode
R14212 N14211 N14212 10
D14212 N14212 0 diode
R14213 N14212 N14213 10
D14213 N14213 0 diode
R14214 N14213 N14214 10
D14214 N14214 0 diode
R14215 N14214 N14215 10
D14215 N14215 0 diode
R14216 N14215 N14216 10
D14216 N14216 0 diode
R14217 N14216 N14217 10
D14217 N14217 0 diode
R14218 N14217 N14218 10
D14218 N14218 0 diode
R14219 N14218 N14219 10
D14219 N14219 0 diode
R14220 N14219 N14220 10
D14220 N14220 0 diode
R14221 N14220 N14221 10
D14221 N14221 0 diode
R14222 N14221 N14222 10
D14222 N14222 0 diode
R14223 N14222 N14223 10
D14223 N14223 0 diode
R14224 N14223 N14224 10
D14224 N14224 0 diode
R14225 N14224 N14225 10
D14225 N14225 0 diode
R14226 N14225 N14226 10
D14226 N14226 0 diode
R14227 N14226 N14227 10
D14227 N14227 0 diode
R14228 N14227 N14228 10
D14228 N14228 0 diode
R14229 N14228 N14229 10
D14229 N14229 0 diode
R14230 N14229 N14230 10
D14230 N14230 0 diode
R14231 N14230 N14231 10
D14231 N14231 0 diode
R14232 N14231 N14232 10
D14232 N14232 0 diode
R14233 N14232 N14233 10
D14233 N14233 0 diode
R14234 N14233 N14234 10
D14234 N14234 0 diode
R14235 N14234 N14235 10
D14235 N14235 0 diode
R14236 N14235 N14236 10
D14236 N14236 0 diode
R14237 N14236 N14237 10
D14237 N14237 0 diode
R14238 N14237 N14238 10
D14238 N14238 0 diode
R14239 N14238 N14239 10
D14239 N14239 0 diode
R14240 N14239 N14240 10
D14240 N14240 0 diode
R14241 N14240 N14241 10
D14241 N14241 0 diode
R14242 N14241 N14242 10
D14242 N14242 0 diode
R14243 N14242 N14243 10
D14243 N14243 0 diode
R14244 N14243 N14244 10
D14244 N14244 0 diode
R14245 N14244 N14245 10
D14245 N14245 0 diode
R14246 N14245 N14246 10
D14246 N14246 0 diode
R14247 N14246 N14247 10
D14247 N14247 0 diode
R14248 N14247 N14248 10
D14248 N14248 0 diode
R14249 N14248 N14249 10
D14249 N14249 0 diode
R14250 N14249 N14250 10
D14250 N14250 0 diode
R14251 N14250 N14251 10
D14251 N14251 0 diode
R14252 N14251 N14252 10
D14252 N14252 0 diode
R14253 N14252 N14253 10
D14253 N14253 0 diode
R14254 N14253 N14254 10
D14254 N14254 0 diode
R14255 N14254 N14255 10
D14255 N14255 0 diode
R14256 N14255 N14256 10
D14256 N14256 0 diode
R14257 N14256 N14257 10
D14257 N14257 0 diode
R14258 N14257 N14258 10
D14258 N14258 0 diode
R14259 N14258 N14259 10
D14259 N14259 0 diode
R14260 N14259 N14260 10
D14260 N14260 0 diode
R14261 N14260 N14261 10
D14261 N14261 0 diode
R14262 N14261 N14262 10
D14262 N14262 0 diode
R14263 N14262 N14263 10
D14263 N14263 0 diode
R14264 N14263 N14264 10
D14264 N14264 0 diode
R14265 N14264 N14265 10
D14265 N14265 0 diode
R14266 N14265 N14266 10
D14266 N14266 0 diode
R14267 N14266 N14267 10
D14267 N14267 0 diode
R14268 N14267 N14268 10
D14268 N14268 0 diode
R14269 N14268 N14269 10
D14269 N14269 0 diode
R14270 N14269 N14270 10
D14270 N14270 0 diode
R14271 N14270 N14271 10
D14271 N14271 0 diode
R14272 N14271 N14272 10
D14272 N14272 0 diode
R14273 N14272 N14273 10
D14273 N14273 0 diode
R14274 N14273 N14274 10
D14274 N14274 0 diode
R14275 N14274 N14275 10
D14275 N14275 0 diode
R14276 N14275 N14276 10
D14276 N14276 0 diode
R14277 N14276 N14277 10
D14277 N14277 0 diode
R14278 N14277 N14278 10
D14278 N14278 0 diode
R14279 N14278 N14279 10
D14279 N14279 0 diode
R14280 N14279 N14280 10
D14280 N14280 0 diode
R14281 N14280 N14281 10
D14281 N14281 0 diode
R14282 N14281 N14282 10
D14282 N14282 0 diode
R14283 N14282 N14283 10
D14283 N14283 0 diode
R14284 N14283 N14284 10
D14284 N14284 0 diode
R14285 N14284 N14285 10
D14285 N14285 0 diode
R14286 N14285 N14286 10
D14286 N14286 0 diode
R14287 N14286 N14287 10
D14287 N14287 0 diode
R14288 N14287 N14288 10
D14288 N14288 0 diode
R14289 N14288 N14289 10
D14289 N14289 0 diode
R14290 N14289 N14290 10
D14290 N14290 0 diode
R14291 N14290 N14291 10
D14291 N14291 0 diode
R14292 N14291 N14292 10
D14292 N14292 0 diode
R14293 N14292 N14293 10
D14293 N14293 0 diode
R14294 N14293 N14294 10
D14294 N14294 0 diode
R14295 N14294 N14295 10
D14295 N14295 0 diode
R14296 N14295 N14296 10
D14296 N14296 0 diode
R14297 N14296 N14297 10
D14297 N14297 0 diode
R14298 N14297 N14298 10
D14298 N14298 0 diode
R14299 N14298 N14299 10
D14299 N14299 0 diode
R14300 N14299 N14300 10
D14300 N14300 0 diode
R14301 N14300 N14301 10
D14301 N14301 0 diode
R14302 N14301 N14302 10
D14302 N14302 0 diode
R14303 N14302 N14303 10
D14303 N14303 0 diode
R14304 N14303 N14304 10
D14304 N14304 0 diode
R14305 N14304 N14305 10
D14305 N14305 0 diode
R14306 N14305 N14306 10
D14306 N14306 0 diode
R14307 N14306 N14307 10
D14307 N14307 0 diode
R14308 N14307 N14308 10
D14308 N14308 0 diode
R14309 N14308 N14309 10
D14309 N14309 0 diode
R14310 N14309 N14310 10
D14310 N14310 0 diode
R14311 N14310 N14311 10
D14311 N14311 0 diode
R14312 N14311 N14312 10
D14312 N14312 0 diode
R14313 N14312 N14313 10
D14313 N14313 0 diode
R14314 N14313 N14314 10
D14314 N14314 0 diode
R14315 N14314 N14315 10
D14315 N14315 0 diode
R14316 N14315 N14316 10
D14316 N14316 0 diode
R14317 N14316 N14317 10
D14317 N14317 0 diode
R14318 N14317 N14318 10
D14318 N14318 0 diode
R14319 N14318 N14319 10
D14319 N14319 0 diode
R14320 N14319 N14320 10
D14320 N14320 0 diode
R14321 N14320 N14321 10
D14321 N14321 0 diode
R14322 N14321 N14322 10
D14322 N14322 0 diode
R14323 N14322 N14323 10
D14323 N14323 0 diode
R14324 N14323 N14324 10
D14324 N14324 0 diode
R14325 N14324 N14325 10
D14325 N14325 0 diode
R14326 N14325 N14326 10
D14326 N14326 0 diode
R14327 N14326 N14327 10
D14327 N14327 0 diode
R14328 N14327 N14328 10
D14328 N14328 0 diode
R14329 N14328 N14329 10
D14329 N14329 0 diode
R14330 N14329 N14330 10
D14330 N14330 0 diode
R14331 N14330 N14331 10
D14331 N14331 0 diode
R14332 N14331 N14332 10
D14332 N14332 0 diode
R14333 N14332 N14333 10
D14333 N14333 0 diode
R14334 N14333 N14334 10
D14334 N14334 0 diode
R14335 N14334 N14335 10
D14335 N14335 0 diode
R14336 N14335 N14336 10
D14336 N14336 0 diode
R14337 N14336 N14337 10
D14337 N14337 0 diode
R14338 N14337 N14338 10
D14338 N14338 0 diode
R14339 N14338 N14339 10
D14339 N14339 0 diode
R14340 N14339 N14340 10
D14340 N14340 0 diode
R14341 N14340 N14341 10
D14341 N14341 0 diode
R14342 N14341 N14342 10
D14342 N14342 0 diode
R14343 N14342 N14343 10
D14343 N14343 0 diode
R14344 N14343 N14344 10
D14344 N14344 0 diode
R14345 N14344 N14345 10
D14345 N14345 0 diode
R14346 N14345 N14346 10
D14346 N14346 0 diode
R14347 N14346 N14347 10
D14347 N14347 0 diode
R14348 N14347 N14348 10
D14348 N14348 0 diode
R14349 N14348 N14349 10
D14349 N14349 0 diode
R14350 N14349 N14350 10
D14350 N14350 0 diode
R14351 N14350 N14351 10
D14351 N14351 0 diode
R14352 N14351 N14352 10
D14352 N14352 0 diode
R14353 N14352 N14353 10
D14353 N14353 0 diode
R14354 N14353 N14354 10
D14354 N14354 0 diode
R14355 N14354 N14355 10
D14355 N14355 0 diode
R14356 N14355 N14356 10
D14356 N14356 0 diode
R14357 N14356 N14357 10
D14357 N14357 0 diode
R14358 N14357 N14358 10
D14358 N14358 0 diode
R14359 N14358 N14359 10
D14359 N14359 0 diode
R14360 N14359 N14360 10
D14360 N14360 0 diode
R14361 N14360 N14361 10
D14361 N14361 0 diode
R14362 N14361 N14362 10
D14362 N14362 0 diode
R14363 N14362 N14363 10
D14363 N14363 0 diode
R14364 N14363 N14364 10
D14364 N14364 0 diode
R14365 N14364 N14365 10
D14365 N14365 0 diode
R14366 N14365 N14366 10
D14366 N14366 0 diode
R14367 N14366 N14367 10
D14367 N14367 0 diode
R14368 N14367 N14368 10
D14368 N14368 0 diode
R14369 N14368 N14369 10
D14369 N14369 0 diode
R14370 N14369 N14370 10
D14370 N14370 0 diode
R14371 N14370 N14371 10
D14371 N14371 0 diode
R14372 N14371 N14372 10
D14372 N14372 0 diode
R14373 N14372 N14373 10
D14373 N14373 0 diode
R14374 N14373 N14374 10
D14374 N14374 0 diode
R14375 N14374 N14375 10
D14375 N14375 0 diode
R14376 N14375 N14376 10
D14376 N14376 0 diode
R14377 N14376 N14377 10
D14377 N14377 0 diode
R14378 N14377 N14378 10
D14378 N14378 0 diode
R14379 N14378 N14379 10
D14379 N14379 0 diode
R14380 N14379 N14380 10
D14380 N14380 0 diode
R14381 N14380 N14381 10
D14381 N14381 0 diode
R14382 N14381 N14382 10
D14382 N14382 0 diode
R14383 N14382 N14383 10
D14383 N14383 0 diode
R14384 N14383 N14384 10
D14384 N14384 0 diode
R14385 N14384 N14385 10
D14385 N14385 0 diode
R14386 N14385 N14386 10
D14386 N14386 0 diode
R14387 N14386 N14387 10
D14387 N14387 0 diode
R14388 N14387 N14388 10
D14388 N14388 0 diode
R14389 N14388 N14389 10
D14389 N14389 0 diode
R14390 N14389 N14390 10
D14390 N14390 0 diode
R14391 N14390 N14391 10
D14391 N14391 0 diode
R14392 N14391 N14392 10
D14392 N14392 0 diode
R14393 N14392 N14393 10
D14393 N14393 0 diode
R14394 N14393 N14394 10
D14394 N14394 0 diode
R14395 N14394 N14395 10
D14395 N14395 0 diode
R14396 N14395 N14396 10
D14396 N14396 0 diode
R14397 N14396 N14397 10
D14397 N14397 0 diode
R14398 N14397 N14398 10
D14398 N14398 0 diode
R14399 N14398 N14399 10
D14399 N14399 0 diode
R14400 N14399 N14400 10
D14400 N14400 0 diode
R14401 N14400 N14401 10
D14401 N14401 0 diode
R14402 N14401 N14402 10
D14402 N14402 0 diode
R14403 N14402 N14403 10
D14403 N14403 0 diode
R14404 N14403 N14404 10
D14404 N14404 0 diode
R14405 N14404 N14405 10
D14405 N14405 0 diode
R14406 N14405 N14406 10
D14406 N14406 0 diode
R14407 N14406 N14407 10
D14407 N14407 0 diode
R14408 N14407 N14408 10
D14408 N14408 0 diode
R14409 N14408 N14409 10
D14409 N14409 0 diode
R14410 N14409 N14410 10
D14410 N14410 0 diode
R14411 N14410 N14411 10
D14411 N14411 0 diode
R14412 N14411 N14412 10
D14412 N14412 0 diode
R14413 N14412 N14413 10
D14413 N14413 0 diode
R14414 N14413 N14414 10
D14414 N14414 0 diode
R14415 N14414 N14415 10
D14415 N14415 0 diode
R14416 N14415 N14416 10
D14416 N14416 0 diode
R14417 N14416 N14417 10
D14417 N14417 0 diode
R14418 N14417 N14418 10
D14418 N14418 0 diode
R14419 N14418 N14419 10
D14419 N14419 0 diode
R14420 N14419 N14420 10
D14420 N14420 0 diode
R14421 N14420 N14421 10
D14421 N14421 0 diode
R14422 N14421 N14422 10
D14422 N14422 0 diode
R14423 N14422 N14423 10
D14423 N14423 0 diode
R14424 N14423 N14424 10
D14424 N14424 0 diode
R14425 N14424 N14425 10
D14425 N14425 0 diode
R14426 N14425 N14426 10
D14426 N14426 0 diode
R14427 N14426 N14427 10
D14427 N14427 0 diode
R14428 N14427 N14428 10
D14428 N14428 0 diode
R14429 N14428 N14429 10
D14429 N14429 0 diode
R14430 N14429 N14430 10
D14430 N14430 0 diode
R14431 N14430 N14431 10
D14431 N14431 0 diode
R14432 N14431 N14432 10
D14432 N14432 0 diode
R14433 N14432 N14433 10
D14433 N14433 0 diode
R14434 N14433 N14434 10
D14434 N14434 0 diode
R14435 N14434 N14435 10
D14435 N14435 0 diode
R14436 N14435 N14436 10
D14436 N14436 0 diode
R14437 N14436 N14437 10
D14437 N14437 0 diode
R14438 N14437 N14438 10
D14438 N14438 0 diode
R14439 N14438 N14439 10
D14439 N14439 0 diode
R14440 N14439 N14440 10
D14440 N14440 0 diode
R14441 N14440 N14441 10
D14441 N14441 0 diode
R14442 N14441 N14442 10
D14442 N14442 0 diode
R14443 N14442 N14443 10
D14443 N14443 0 diode
R14444 N14443 N14444 10
D14444 N14444 0 diode
R14445 N14444 N14445 10
D14445 N14445 0 diode
R14446 N14445 N14446 10
D14446 N14446 0 diode
R14447 N14446 N14447 10
D14447 N14447 0 diode
R14448 N14447 N14448 10
D14448 N14448 0 diode
R14449 N14448 N14449 10
D14449 N14449 0 diode
R14450 N14449 N14450 10
D14450 N14450 0 diode
R14451 N14450 N14451 10
D14451 N14451 0 diode
R14452 N14451 N14452 10
D14452 N14452 0 diode
R14453 N14452 N14453 10
D14453 N14453 0 diode
R14454 N14453 N14454 10
D14454 N14454 0 diode
R14455 N14454 N14455 10
D14455 N14455 0 diode
R14456 N14455 N14456 10
D14456 N14456 0 diode
R14457 N14456 N14457 10
D14457 N14457 0 diode
R14458 N14457 N14458 10
D14458 N14458 0 diode
R14459 N14458 N14459 10
D14459 N14459 0 diode
R14460 N14459 N14460 10
D14460 N14460 0 diode
R14461 N14460 N14461 10
D14461 N14461 0 diode
R14462 N14461 N14462 10
D14462 N14462 0 diode
R14463 N14462 N14463 10
D14463 N14463 0 diode
R14464 N14463 N14464 10
D14464 N14464 0 diode
R14465 N14464 N14465 10
D14465 N14465 0 diode
R14466 N14465 N14466 10
D14466 N14466 0 diode
R14467 N14466 N14467 10
D14467 N14467 0 diode
R14468 N14467 N14468 10
D14468 N14468 0 diode
R14469 N14468 N14469 10
D14469 N14469 0 diode
R14470 N14469 N14470 10
D14470 N14470 0 diode
R14471 N14470 N14471 10
D14471 N14471 0 diode
R14472 N14471 N14472 10
D14472 N14472 0 diode
R14473 N14472 N14473 10
D14473 N14473 0 diode
R14474 N14473 N14474 10
D14474 N14474 0 diode
R14475 N14474 N14475 10
D14475 N14475 0 diode
R14476 N14475 N14476 10
D14476 N14476 0 diode
R14477 N14476 N14477 10
D14477 N14477 0 diode
R14478 N14477 N14478 10
D14478 N14478 0 diode
R14479 N14478 N14479 10
D14479 N14479 0 diode
R14480 N14479 N14480 10
D14480 N14480 0 diode
R14481 N14480 N14481 10
D14481 N14481 0 diode
R14482 N14481 N14482 10
D14482 N14482 0 diode
R14483 N14482 N14483 10
D14483 N14483 0 diode
R14484 N14483 N14484 10
D14484 N14484 0 diode
R14485 N14484 N14485 10
D14485 N14485 0 diode
R14486 N14485 N14486 10
D14486 N14486 0 diode
R14487 N14486 N14487 10
D14487 N14487 0 diode
R14488 N14487 N14488 10
D14488 N14488 0 diode
R14489 N14488 N14489 10
D14489 N14489 0 diode
R14490 N14489 N14490 10
D14490 N14490 0 diode
R14491 N14490 N14491 10
D14491 N14491 0 diode
R14492 N14491 N14492 10
D14492 N14492 0 diode
R14493 N14492 N14493 10
D14493 N14493 0 diode
R14494 N14493 N14494 10
D14494 N14494 0 diode
R14495 N14494 N14495 10
D14495 N14495 0 diode
R14496 N14495 N14496 10
D14496 N14496 0 diode
R14497 N14496 N14497 10
D14497 N14497 0 diode
R14498 N14497 N14498 10
D14498 N14498 0 diode
R14499 N14498 N14499 10
D14499 N14499 0 diode
R14500 N14499 N14500 10
D14500 N14500 0 diode
R14501 N14500 N14501 10
D14501 N14501 0 diode
R14502 N14501 N14502 10
D14502 N14502 0 diode
R14503 N14502 N14503 10
D14503 N14503 0 diode
R14504 N14503 N14504 10
D14504 N14504 0 diode
R14505 N14504 N14505 10
D14505 N14505 0 diode
R14506 N14505 N14506 10
D14506 N14506 0 diode
R14507 N14506 N14507 10
D14507 N14507 0 diode
R14508 N14507 N14508 10
D14508 N14508 0 diode
R14509 N14508 N14509 10
D14509 N14509 0 diode
R14510 N14509 N14510 10
D14510 N14510 0 diode
R14511 N14510 N14511 10
D14511 N14511 0 diode
R14512 N14511 N14512 10
D14512 N14512 0 diode
R14513 N14512 N14513 10
D14513 N14513 0 diode
R14514 N14513 N14514 10
D14514 N14514 0 diode
R14515 N14514 N14515 10
D14515 N14515 0 diode
R14516 N14515 N14516 10
D14516 N14516 0 diode
R14517 N14516 N14517 10
D14517 N14517 0 diode
R14518 N14517 N14518 10
D14518 N14518 0 diode
R14519 N14518 N14519 10
D14519 N14519 0 diode
R14520 N14519 N14520 10
D14520 N14520 0 diode
R14521 N14520 N14521 10
D14521 N14521 0 diode
R14522 N14521 N14522 10
D14522 N14522 0 diode
R14523 N14522 N14523 10
D14523 N14523 0 diode
R14524 N14523 N14524 10
D14524 N14524 0 diode
R14525 N14524 N14525 10
D14525 N14525 0 diode
R14526 N14525 N14526 10
D14526 N14526 0 diode
R14527 N14526 N14527 10
D14527 N14527 0 diode
R14528 N14527 N14528 10
D14528 N14528 0 diode
R14529 N14528 N14529 10
D14529 N14529 0 diode
R14530 N14529 N14530 10
D14530 N14530 0 diode
R14531 N14530 N14531 10
D14531 N14531 0 diode
R14532 N14531 N14532 10
D14532 N14532 0 diode
R14533 N14532 N14533 10
D14533 N14533 0 diode
R14534 N14533 N14534 10
D14534 N14534 0 diode
R14535 N14534 N14535 10
D14535 N14535 0 diode
R14536 N14535 N14536 10
D14536 N14536 0 diode
R14537 N14536 N14537 10
D14537 N14537 0 diode
R14538 N14537 N14538 10
D14538 N14538 0 diode
R14539 N14538 N14539 10
D14539 N14539 0 diode
R14540 N14539 N14540 10
D14540 N14540 0 diode
R14541 N14540 N14541 10
D14541 N14541 0 diode
R14542 N14541 N14542 10
D14542 N14542 0 diode
R14543 N14542 N14543 10
D14543 N14543 0 diode
R14544 N14543 N14544 10
D14544 N14544 0 diode
R14545 N14544 N14545 10
D14545 N14545 0 diode
R14546 N14545 N14546 10
D14546 N14546 0 diode
R14547 N14546 N14547 10
D14547 N14547 0 diode
R14548 N14547 N14548 10
D14548 N14548 0 diode
R14549 N14548 N14549 10
D14549 N14549 0 diode
R14550 N14549 N14550 10
D14550 N14550 0 diode
R14551 N14550 N14551 10
D14551 N14551 0 diode
R14552 N14551 N14552 10
D14552 N14552 0 diode
R14553 N14552 N14553 10
D14553 N14553 0 diode
R14554 N14553 N14554 10
D14554 N14554 0 diode
R14555 N14554 N14555 10
D14555 N14555 0 diode
R14556 N14555 N14556 10
D14556 N14556 0 diode
R14557 N14556 N14557 10
D14557 N14557 0 diode
R14558 N14557 N14558 10
D14558 N14558 0 diode
R14559 N14558 N14559 10
D14559 N14559 0 diode
R14560 N14559 N14560 10
D14560 N14560 0 diode
R14561 N14560 N14561 10
D14561 N14561 0 diode
R14562 N14561 N14562 10
D14562 N14562 0 diode
R14563 N14562 N14563 10
D14563 N14563 0 diode
R14564 N14563 N14564 10
D14564 N14564 0 diode
R14565 N14564 N14565 10
D14565 N14565 0 diode
R14566 N14565 N14566 10
D14566 N14566 0 diode
R14567 N14566 N14567 10
D14567 N14567 0 diode
R14568 N14567 N14568 10
D14568 N14568 0 diode
R14569 N14568 N14569 10
D14569 N14569 0 diode
R14570 N14569 N14570 10
D14570 N14570 0 diode
R14571 N14570 N14571 10
D14571 N14571 0 diode
R14572 N14571 N14572 10
D14572 N14572 0 diode
R14573 N14572 N14573 10
D14573 N14573 0 diode
R14574 N14573 N14574 10
D14574 N14574 0 diode
R14575 N14574 N14575 10
D14575 N14575 0 diode
R14576 N14575 N14576 10
D14576 N14576 0 diode
R14577 N14576 N14577 10
D14577 N14577 0 diode
R14578 N14577 N14578 10
D14578 N14578 0 diode
R14579 N14578 N14579 10
D14579 N14579 0 diode
R14580 N14579 N14580 10
D14580 N14580 0 diode
R14581 N14580 N14581 10
D14581 N14581 0 diode
R14582 N14581 N14582 10
D14582 N14582 0 diode
R14583 N14582 N14583 10
D14583 N14583 0 diode
R14584 N14583 N14584 10
D14584 N14584 0 diode
R14585 N14584 N14585 10
D14585 N14585 0 diode
R14586 N14585 N14586 10
D14586 N14586 0 diode
R14587 N14586 N14587 10
D14587 N14587 0 diode
R14588 N14587 N14588 10
D14588 N14588 0 diode
R14589 N14588 N14589 10
D14589 N14589 0 diode
R14590 N14589 N14590 10
D14590 N14590 0 diode
R14591 N14590 N14591 10
D14591 N14591 0 diode
R14592 N14591 N14592 10
D14592 N14592 0 diode
R14593 N14592 N14593 10
D14593 N14593 0 diode
R14594 N14593 N14594 10
D14594 N14594 0 diode
R14595 N14594 N14595 10
D14595 N14595 0 diode
R14596 N14595 N14596 10
D14596 N14596 0 diode
R14597 N14596 N14597 10
D14597 N14597 0 diode
R14598 N14597 N14598 10
D14598 N14598 0 diode
R14599 N14598 N14599 10
D14599 N14599 0 diode
R14600 N14599 N14600 10
D14600 N14600 0 diode
R14601 N14600 N14601 10
D14601 N14601 0 diode
R14602 N14601 N14602 10
D14602 N14602 0 diode
R14603 N14602 N14603 10
D14603 N14603 0 diode
R14604 N14603 N14604 10
D14604 N14604 0 diode
R14605 N14604 N14605 10
D14605 N14605 0 diode
R14606 N14605 N14606 10
D14606 N14606 0 diode
R14607 N14606 N14607 10
D14607 N14607 0 diode
R14608 N14607 N14608 10
D14608 N14608 0 diode
R14609 N14608 N14609 10
D14609 N14609 0 diode
R14610 N14609 N14610 10
D14610 N14610 0 diode
R14611 N14610 N14611 10
D14611 N14611 0 diode
R14612 N14611 N14612 10
D14612 N14612 0 diode
R14613 N14612 N14613 10
D14613 N14613 0 diode
R14614 N14613 N14614 10
D14614 N14614 0 diode
R14615 N14614 N14615 10
D14615 N14615 0 diode
R14616 N14615 N14616 10
D14616 N14616 0 diode
R14617 N14616 N14617 10
D14617 N14617 0 diode
R14618 N14617 N14618 10
D14618 N14618 0 diode
R14619 N14618 N14619 10
D14619 N14619 0 diode
R14620 N14619 N14620 10
D14620 N14620 0 diode
R14621 N14620 N14621 10
D14621 N14621 0 diode
R14622 N14621 N14622 10
D14622 N14622 0 diode
R14623 N14622 N14623 10
D14623 N14623 0 diode
R14624 N14623 N14624 10
D14624 N14624 0 diode
R14625 N14624 N14625 10
D14625 N14625 0 diode
R14626 N14625 N14626 10
D14626 N14626 0 diode
R14627 N14626 N14627 10
D14627 N14627 0 diode
R14628 N14627 N14628 10
D14628 N14628 0 diode
R14629 N14628 N14629 10
D14629 N14629 0 diode
R14630 N14629 N14630 10
D14630 N14630 0 diode
R14631 N14630 N14631 10
D14631 N14631 0 diode
R14632 N14631 N14632 10
D14632 N14632 0 diode
R14633 N14632 N14633 10
D14633 N14633 0 diode
R14634 N14633 N14634 10
D14634 N14634 0 diode
R14635 N14634 N14635 10
D14635 N14635 0 diode
R14636 N14635 N14636 10
D14636 N14636 0 diode
R14637 N14636 N14637 10
D14637 N14637 0 diode
R14638 N14637 N14638 10
D14638 N14638 0 diode
R14639 N14638 N14639 10
D14639 N14639 0 diode
R14640 N14639 N14640 10
D14640 N14640 0 diode
R14641 N14640 N14641 10
D14641 N14641 0 diode
R14642 N14641 N14642 10
D14642 N14642 0 diode
R14643 N14642 N14643 10
D14643 N14643 0 diode
R14644 N14643 N14644 10
D14644 N14644 0 diode
R14645 N14644 N14645 10
D14645 N14645 0 diode
R14646 N14645 N14646 10
D14646 N14646 0 diode
R14647 N14646 N14647 10
D14647 N14647 0 diode
R14648 N14647 N14648 10
D14648 N14648 0 diode
R14649 N14648 N14649 10
D14649 N14649 0 diode
R14650 N14649 N14650 10
D14650 N14650 0 diode
R14651 N14650 N14651 10
D14651 N14651 0 diode
R14652 N14651 N14652 10
D14652 N14652 0 diode
R14653 N14652 N14653 10
D14653 N14653 0 diode
R14654 N14653 N14654 10
D14654 N14654 0 diode
R14655 N14654 N14655 10
D14655 N14655 0 diode
R14656 N14655 N14656 10
D14656 N14656 0 diode
R14657 N14656 N14657 10
D14657 N14657 0 diode
R14658 N14657 N14658 10
D14658 N14658 0 diode
R14659 N14658 N14659 10
D14659 N14659 0 diode
R14660 N14659 N14660 10
D14660 N14660 0 diode
R14661 N14660 N14661 10
D14661 N14661 0 diode
R14662 N14661 N14662 10
D14662 N14662 0 diode
R14663 N14662 N14663 10
D14663 N14663 0 diode
R14664 N14663 N14664 10
D14664 N14664 0 diode
R14665 N14664 N14665 10
D14665 N14665 0 diode
R14666 N14665 N14666 10
D14666 N14666 0 diode
R14667 N14666 N14667 10
D14667 N14667 0 diode
R14668 N14667 N14668 10
D14668 N14668 0 diode
R14669 N14668 N14669 10
D14669 N14669 0 diode
R14670 N14669 N14670 10
D14670 N14670 0 diode
R14671 N14670 N14671 10
D14671 N14671 0 diode
R14672 N14671 N14672 10
D14672 N14672 0 diode
R14673 N14672 N14673 10
D14673 N14673 0 diode
R14674 N14673 N14674 10
D14674 N14674 0 diode
R14675 N14674 N14675 10
D14675 N14675 0 diode
R14676 N14675 N14676 10
D14676 N14676 0 diode
R14677 N14676 N14677 10
D14677 N14677 0 diode
R14678 N14677 N14678 10
D14678 N14678 0 diode
R14679 N14678 N14679 10
D14679 N14679 0 diode
R14680 N14679 N14680 10
D14680 N14680 0 diode
R14681 N14680 N14681 10
D14681 N14681 0 diode
R14682 N14681 N14682 10
D14682 N14682 0 diode
R14683 N14682 N14683 10
D14683 N14683 0 diode
R14684 N14683 N14684 10
D14684 N14684 0 diode
R14685 N14684 N14685 10
D14685 N14685 0 diode
R14686 N14685 N14686 10
D14686 N14686 0 diode
R14687 N14686 N14687 10
D14687 N14687 0 diode
R14688 N14687 N14688 10
D14688 N14688 0 diode
R14689 N14688 N14689 10
D14689 N14689 0 diode
R14690 N14689 N14690 10
D14690 N14690 0 diode
R14691 N14690 N14691 10
D14691 N14691 0 diode
R14692 N14691 N14692 10
D14692 N14692 0 diode
R14693 N14692 N14693 10
D14693 N14693 0 diode
R14694 N14693 N14694 10
D14694 N14694 0 diode
R14695 N14694 N14695 10
D14695 N14695 0 diode
R14696 N14695 N14696 10
D14696 N14696 0 diode
R14697 N14696 N14697 10
D14697 N14697 0 diode
R14698 N14697 N14698 10
D14698 N14698 0 diode
R14699 N14698 N14699 10
D14699 N14699 0 diode
R14700 N14699 N14700 10
D14700 N14700 0 diode
R14701 N14700 N14701 10
D14701 N14701 0 diode
R14702 N14701 N14702 10
D14702 N14702 0 diode
R14703 N14702 N14703 10
D14703 N14703 0 diode
R14704 N14703 N14704 10
D14704 N14704 0 diode
R14705 N14704 N14705 10
D14705 N14705 0 diode
R14706 N14705 N14706 10
D14706 N14706 0 diode
R14707 N14706 N14707 10
D14707 N14707 0 diode
R14708 N14707 N14708 10
D14708 N14708 0 diode
R14709 N14708 N14709 10
D14709 N14709 0 diode
R14710 N14709 N14710 10
D14710 N14710 0 diode
R14711 N14710 N14711 10
D14711 N14711 0 diode
R14712 N14711 N14712 10
D14712 N14712 0 diode
R14713 N14712 N14713 10
D14713 N14713 0 diode
R14714 N14713 N14714 10
D14714 N14714 0 diode
R14715 N14714 N14715 10
D14715 N14715 0 diode
R14716 N14715 N14716 10
D14716 N14716 0 diode
R14717 N14716 N14717 10
D14717 N14717 0 diode
R14718 N14717 N14718 10
D14718 N14718 0 diode
R14719 N14718 N14719 10
D14719 N14719 0 diode
R14720 N14719 N14720 10
D14720 N14720 0 diode
R14721 N14720 N14721 10
D14721 N14721 0 diode
R14722 N14721 N14722 10
D14722 N14722 0 diode
R14723 N14722 N14723 10
D14723 N14723 0 diode
R14724 N14723 N14724 10
D14724 N14724 0 diode
R14725 N14724 N14725 10
D14725 N14725 0 diode
R14726 N14725 N14726 10
D14726 N14726 0 diode
R14727 N14726 N14727 10
D14727 N14727 0 diode
R14728 N14727 N14728 10
D14728 N14728 0 diode
R14729 N14728 N14729 10
D14729 N14729 0 diode
R14730 N14729 N14730 10
D14730 N14730 0 diode
R14731 N14730 N14731 10
D14731 N14731 0 diode
R14732 N14731 N14732 10
D14732 N14732 0 diode
R14733 N14732 N14733 10
D14733 N14733 0 diode
R14734 N14733 N14734 10
D14734 N14734 0 diode
R14735 N14734 N14735 10
D14735 N14735 0 diode
R14736 N14735 N14736 10
D14736 N14736 0 diode
R14737 N14736 N14737 10
D14737 N14737 0 diode
R14738 N14737 N14738 10
D14738 N14738 0 diode
R14739 N14738 N14739 10
D14739 N14739 0 diode
R14740 N14739 N14740 10
D14740 N14740 0 diode
R14741 N14740 N14741 10
D14741 N14741 0 diode
R14742 N14741 N14742 10
D14742 N14742 0 diode
R14743 N14742 N14743 10
D14743 N14743 0 diode
R14744 N14743 N14744 10
D14744 N14744 0 diode
R14745 N14744 N14745 10
D14745 N14745 0 diode
R14746 N14745 N14746 10
D14746 N14746 0 diode
R14747 N14746 N14747 10
D14747 N14747 0 diode
R14748 N14747 N14748 10
D14748 N14748 0 diode
R14749 N14748 N14749 10
D14749 N14749 0 diode
R14750 N14749 N14750 10
D14750 N14750 0 diode
R14751 N14750 N14751 10
D14751 N14751 0 diode
R14752 N14751 N14752 10
D14752 N14752 0 diode
R14753 N14752 N14753 10
D14753 N14753 0 diode
R14754 N14753 N14754 10
D14754 N14754 0 diode
R14755 N14754 N14755 10
D14755 N14755 0 diode
R14756 N14755 N14756 10
D14756 N14756 0 diode
R14757 N14756 N14757 10
D14757 N14757 0 diode
R14758 N14757 N14758 10
D14758 N14758 0 diode
R14759 N14758 N14759 10
D14759 N14759 0 diode
R14760 N14759 N14760 10
D14760 N14760 0 diode
R14761 N14760 N14761 10
D14761 N14761 0 diode
R14762 N14761 N14762 10
D14762 N14762 0 diode
R14763 N14762 N14763 10
D14763 N14763 0 diode
R14764 N14763 N14764 10
D14764 N14764 0 diode
R14765 N14764 N14765 10
D14765 N14765 0 diode
R14766 N14765 N14766 10
D14766 N14766 0 diode
R14767 N14766 N14767 10
D14767 N14767 0 diode
R14768 N14767 N14768 10
D14768 N14768 0 diode
R14769 N14768 N14769 10
D14769 N14769 0 diode
R14770 N14769 N14770 10
D14770 N14770 0 diode
R14771 N14770 N14771 10
D14771 N14771 0 diode
R14772 N14771 N14772 10
D14772 N14772 0 diode
R14773 N14772 N14773 10
D14773 N14773 0 diode
R14774 N14773 N14774 10
D14774 N14774 0 diode
R14775 N14774 N14775 10
D14775 N14775 0 diode
R14776 N14775 N14776 10
D14776 N14776 0 diode
R14777 N14776 N14777 10
D14777 N14777 0 diode
R14778 N14777 N14778 10
D14778 N14778 0 diode
R14779 N14778 N14779 10
D14779 N14779 0 diode
R14780 N14779 N14780 10
D14780 N14780 0 diode
R14781 N14780 N14781 10
D14781 N14781 0 diode
R14782 N14781 N14782 10
D14782 N14782 0 diode
R14783 N14782 N14783 10
D14783 N14783 0 diode
R14784 N14783 N14784 10
D14784 N14784 0 diode
R14785 N14784 N14785 10
D14785 N14785 0 diode
R14786 N14785 N14786 10
D14786 N14786 0 diode
R14787 N14786 N14787 10
D14787 N14787 0 diode
R14788 N14787 N14788 10
D14788 N14788 0 diode
R14789 N14788 N14789 10
D14789 N14789 0 diode
R14790 N14789 N14790 10
D14790 N14790 0 diode
R14791 N14790 N14791 10
D14791 N14791 0 diode
R14792 N14791 N14792 10
D14792 N14792 0 diode
R14793 N14792 N14793 10
D14793 N14793 0 diode
R14794 N14793 N14794 10
D14794 N14794 0 diode
R14795 N14794 N14795 10
D14795 N14795 0 diode
R14796 N14795 N14796 10
D14796 N14796 0 diode
R14797 N14796 N14797 10
D14797 N14797 0 diode
R14798 N14797 N14798 10
D14798 N14798 0 diode
R14799 N14798 N14799 10
D14799 N14799 0 diode
R14800 N14799 N14800 10
D14800 N14800 0 diode
R14801 N14800 N14801 10
D14801 N14801 0 diode
R14802 N14801 N14802 10
D14802 N14802 0 diode
R14803 N14802 N14803 10
D14803 N14803 0 diode
R14804 N14803 N14804 10
D14804 N14804 0 diode
R14805 N14804 N14805 10
D14805 N14805 0 diode
R14806 N14805 N14806 10
D14806 N14806 0 diode
R14807 N14806 N14807 10
D14807 N14807 0 diode
R14808 N14807 N14808 10
D14808 N14808 0 diode
R14809 N14808 N14809 10
D14809 N14809 0 diode
R14810 N14809 N14810 10
D14810 N14810 0 diode
R14811 N14810 N14811 10
D14811 N14811 0 diode
R14812 N14811 N14812 10
D14812 N14812 0 diode
R14813 N14812 N14813 10
D14813 N14813 0 diode
R14814 N14813 N14814 10
D14814 N14814 0 diode
R14815 N14814 N14815 10
D14815 N14815 0 diode
R14816 N14815 N14816 10
D14816 N14816 0 diode
R14817 N14816 N14817 10
D14817 N14817 0 diode
R14818 N14817 N14818 10
D14818 N14818 0 diode
R14819 N14818 N14819 10
D14819 N14819 0 diode
R14820 N14819 N14820 10
D14820 N14820 0 diode
R14821 N14820 N14821 10
D14821 N14821 0 diode
R14822 N14821 N14822 10
D14822 N14822 0 diode
R14823 N14822 N14823 10
D14823 N14823 0 diode
R14824 N14823 N14824 10
D14824 N14824 0 diode
R14825 N14824 N14825 10
D14825 N14825 0 diode
R14826 N14825 N14826 10
D14826 N14826 0 diode
R14827 N14826 N14827 10
D14827 N14827 0 diode
R14828 N14827 N14828 10
D14828 N14828 0 diode
R14829 N14828 N14829 10
D14829 N14829 0 diode
R14830 N14829 N14830 10
D14830 N14830 0 diode
R14831 N14830 N14831 10
D14831 N14831 0 diode
R14832 N14831 N14832 10
D14832 N14832 0 diode
R14833 N14832 N14833 10
D14833 N14833 0 diode
R14834 N14833 N14834 10
D14834 N14834 0 diode
R14835 N14834 N14835 10
D14835 N14835 0 diode
R14836 N14835 N14836 10
D14836 N14836 0 diode
R14837 N14836 N14837 10
D14837 N14837 0 diode
R14838 N14837 N14838 10
D14838 N14838 0 diode
R14839 N14838 N14839 10
D14839 N14839 0 diode
R14840 N14839 N14840 10
D14840 N14840 0 diode
R14841 N14840 N14841 10
D14841 N14841 0 diode
R14842 N14841 N14842 10
D14842 N14842 0 diode
R14843 N14842 N14843 10
D14843 N14843 0 diode
R14844 N14843 N14844 10
D14844 N14844 0 diode
R14845 N14844 N14845 10
D14845 N14845 0 diode
R14846 N14845 N14846 10
D14846 N14846 0 diode
R14847 N14846 N14847 10
D14847 N14847 0 diode
R14848 N14847 N14848 10
D14848 N14848 0 diode
R14849 N14848 N14849 10
D14849 N14849 0 diode
R14850 N14849 N14850 10
D14850 N14850 0 diode
R14851 N14850 N14851 10
D14851 N14851 0 diode
R14852 N14851 N14852 10
D14852 N14852 0 diode
R14853 N14852 N14853 10
D14853 N14853 0 diode
R14854 N14853 N14854 10
D14854 N14854 0 diode
R14855 N14854 N14855 10
D14855 N14855 0 diode
R14856 N14855 N14856 10
D14856 N14856 0 diode
R14857 N14856 N14857 10
D14857 N14857 0 diode
R14858 N14857 N14858 10
D14858 N14858 0 diode
R14859 N14858 N14859 10
D14859 N14859 0 diode
R14860 N14859 N14860 10
D14860 N14860 0 diode
R14861 N14860 N14861 10
D14861 N14861 0 diode
R14862 N14861 N14862 10
D14862 N14862 0 diode
R14863 N14862 N14863 10
D14863 N14863 0 diode
R14864 N14863 N14864 10
D14864 N14864 0 diode
R14865 N14864 N14865 10
D14865 N14865 0 diode
R14866 N14865 N14866 10
D14866 N14866 0 diode
R14867 N14866 N14867 10
D14867 N14867 0 diode
R14868 N14867 N14868 10
D14868 N14868 0 diode
R14869 N14868 N14869 10
D14869 N14869 0 diode
R14870 N14869 N14870 10
D14870 N14870 0 diode
R14871 N14870 N14871 10
D14871 N14871 0 diode
R14872 N14871 N14872 10
D14872 N14872 0 diode
R14873 N14872 N14873 10
D14873 N14873 0 diode
R14874 N14873 N14874 10
D14874 N14874 0 diode
R14875 N14874 N14875 10
D14875 N14875 0 diode
R14876 N14875 N14876 10
D14876 N14876 0 diode
R14877 N14876 N14877 10
D14877 N14877 0 diode
R14878 N14877 N14878 10
D14878 N14878 0 diode
R14879 N14878 N14879 10
D14879 N14879 0 diode
R14880 N14879 N14880 10
D14880 N14880 0 diode
R14881 N14880 N14881 10
D14881 N14881 0 diode
R14882 N14881 N14882 10
D14882 N14882 0 diode
R14883 N14882 N14883 10
D14883 N14883 0 diode
R14884 N14883 N14884 10
D14884 N14884 0 diode
R14885 N14884 N14885 10
D14885 N14885 0 diode
R14886 N14885 N14886 10
D14886 N14886 0 diode
R14887 N14886 N14887 10
D14887 N14887 0 diode
R14888 N14887 N14888 10
D14888 N14888 0 diode
R14889 N14888 N14889 10
D14889 N14889 0 diode
R14890 N14889 N14890 10
D14890 N14890 0 diode
R14891 N14890 N14891 10
D14891 N14891 0 diode
R14892 N14891 N14892 10
D14892 N14892 0 diode
R14893 N14892 N14893 10
D14893 N14893 0 diode
R14894 N14893 N14894 10
D14894 N14894 0 diode
R14895 N14894 N14895 10
D14895 N14895 0 diode
R14896 N14895 N14896 10
D14896 N14896 0 diode
R14897 N14896 N14897 10
D14897 N14897 0 diode
R14898 N14897 N14898 10
D14898 N14898 0 diode
R14899 N14898 N14899 10
D14899 N14899 0 diode
R14900 N14899 N14900 10
D14900 N14900 0 diode
R14901 N14900 N14901 10
D14901 N14901 0 diode
R14902 N14901 N14902 10
D14902 N14902 0 diode
R14903 N14902 N14903 10
D14903 N14903 0 diode
R14904 N14903 N14904 10
D14904 N14904 0 diode
R14905 N14904 N14905 10
D14905 N14905 0 diode
R14906 N14905 N14906 10
D14906 N14906 0 diode
R14907 N14906 N14907 10
D14907 N14907 0 diode
R14908 N14907 N14908 10
D14908 N14908 0 diode
R14909 N14908 N14909 10
D14909 N14909 0 diode
R14910 N14909 N14910 10
D14910 N14910 0 diode
R14911 N14910 N14911 10
D14911 N14911 0 diode
R14912 N14911 N14912 10
D14912 N14912 0 diode
R14913 N14912 N14913 10
D14913 N14913 0 diode
R14914 N14913 N14914 10
D14914 N14914 0 diode
R14915 N14914 N14915 10
D14915 N14915 0 diode
R14916 N14915 N14916 10
D14916 N14916 0 diode
R14917 N14916 N14917 10
D14917 N14917 0 diode
R14918 N14917 N14918 10
D14918 N14918 0 diode
R14919 N14918 N14919 10
D14919 N14919 0 diode
R14920 N14919 N14920 10
D14920 N14920 0 diode
R14921 N14920 N14921 10
D14921 N14921 0 diode
R14922 N14921 N14922 10
D14922 N14922 0 diode
R14923 N14922 N14923 10
D14923 N14923 0 diode
R14924 N14923 N14924 10
D14924 N14924 0 diode
R14925 N14924 N14925 10
D14925 N14925 0 diode
R14926 N14925 N14926 10
D14926 N14926 0 diode
R14927 N14926 N14927 10
D14927 N14927 0 diode
R14928 N14927 N14928 10
D14928 N14928 0 diode
R14929 N14928 N14929 10
D14929 N14929 0 diode
R14930 N14929 N14930 10
D14930 N14930 0 diode
R14931 N14930 N14931 10
D14931 N14931 0 diode
R14932 N14931 N14932 10
D14932 N14932 0 diode
R14933 N14932 N14933 10
D14933 N14933 0 diode
R14934 N14933 N14934 10
D14934 N14934 0 diode
R14935 N14934 N14935 10
D14935 N14935 0 diode
R14936 N14935 N14936 10
D14936 N14936 0 diode
R14937 N14936 N14937 10
D14937 N14937 0 diode
R14938 N14937 N14938 10
D14938 N14938 0 diode
R14939 N14938 N14939 10
D14939 N14939 0 diode
R14940 N14939 N14940 10
D14940 N14940 0 diode
R14941 N14940 N14941 10
D14941 N14941 0 diode
R14942 N14941 N14942 10
D14942 N14942 0 diode
R14943 N14942 N14943 10
D14943 N14943 0 diode
R14944 N14943 N14944 10
D14944 N14944 0 diode
R14945 N14944 N14945 10
D14945 N14945 0 diode
R14946 N14945 N14946 10
D14946 N14946 0 diode
R14947 N14946 N14947 10
D14947 N14947 0 diode
R14948 N14947 N14948 10
D14948 N14948 0 diode
R14949 N14948 N14949 10
D14949 N14949 0 diode
R14950 N14949 N14950 10
D14950 N14950 0 diode
R14951 N14950 N14951 10
D14951 N14951 0 diode
R14952 N14951 N14952 10
D14952 N14952 0 diode
R14953 N14952 N14953 10
D14953 N14953 0 diode
R14954 N14953 N14954 10
D14954 N14954 0 diode
R14955 N14954 N14955 10
D14955 N14955 0 diode
R14956 N14955 N14956 10
D14956 N14956 0 diode
R14957 N14956 N14957 10
D14957 N14957 0 diode
R14958 N14957 N14958 10
D14958 N14958 0 diode
R14959 N14958 N14959 10
D14959 N14959 0 diode
R14960 N14959 N14960 10
D14960 N14960 0 diode
R14961 N14960 N14961 10
D14961 N14961 0 diode
R14962 N14961 N14962 10
D14962 N14962 0 diode
R14963 N14962 N14963 10
D14963 N14963 0 diode
R14964 N14963 N14964 10
D14964 N14964 0 diode
R14965 N14964 N14965 10
D14965 N14965 0 diode
R14966 N14965 N14966 10
D14966 N14966 0 diode
R14967 N14966 N14967 10
D14967 N14967 0 diode
R14968 N14967 N14968 10
D14968 N14968 0 diode
R14969 N14968 N14969 10
D14969 N14969 0 diode
R14970 N14969 N14970 10
D14970 N14970 0 diode
R14971 N14970 N14971 10
D14971 N14971 0 diode
R14972 N14971 N14972 10
D14972 N14972 0 diode
R14973 N14972 N14973 10
D14973 N14973 0 diode
R14974 N14973 N14974 10
D14974 N14974 0 diode
R14975 N14974 N14975 10
D14975 N14975 0 diode
R14976 N14975 N14976 10
D14976 N14976 0 diode
R14977 N14976 N14977 10
D14977 N14977 0 diode
R14978 N14977 N14978 10
D14978 N14978 0 diode
R14979 N14978 N14979 10
D14979 N14979 0 diode
R14980 N14979 N14980 10
D14980 N14980 0 diode
R14981 N14980 N14981 10
D14981 N14981 0 diode
R14982 N14981 N14982 10
D14982 N14982 0 diode
R14983 N14982 N14983 10
D14983 N14983 0 diode
R14984 N14983 N14984 10
D14984 N14984 0 diode
R14985 N14984 N14985 10
D14985 N14985 0 diode
R14986 N14985 N14986 10
D14986 N14986 0 diode
R14987 N14986 N14987 10
D14987 N14987 0 diode
R14988 N14987 N14988 10
D14988 N14988 0 diode
R14989 N14988 N14989 10
D14989 N14989 0 diode
R14990 N14989 N14990 10
D14990 N14990 0 diode
R14991 N14990 N14991 10
D14991 N14991 0 diode
R14992 N14991 N14992 10
D14992 N14992 0 diode
R14993 N14992 N14993 10
D14993 N14993 0 diode
R14994 N14993 N14994 10
D14994 N14994 0 diode
R14995 N14994 N14995 10
D14995 N14995 0 diode
R14996 N14995 N14996 10
D14996 N14996 0 diode
R14997 N14996 N14997 10
D14997 N14997 0 diode
R14998 N14997 N14998 10
D14998 N14998 0 diode
R14999 N14998 N14999 10
D14999 N14999 0 diode
R15000 N14999 N15000 10
D15000 N15000 0 diode
R15001 N15000 N15001 10
D15001 N15001 0 diode
R15002 N15001 N15002 10
D15002 N15002 0 diode
R15003 N15002 N15003 10
D15003 N15003 0 diode
R15004 N15003 N15004 10
D15004 N15004 0 diode
R15005 N15004 N15005 10
D15005 N15005 0 diode
R15006 N15005 N15006 10
D15006 N15006 0 diode
R15007 N15006 N15007 10
D15007 N15007 0 diode
R15008 N15007 N15008 10
D15008 N15008 0 diode
R15009 N15008 N15009 10
D15009 N15009 0 diode
R15010 N15009 N15010 10
D15010 N15010 0 diode
R15011 N15010 N15011 10
D15011 N15011 0 diode
R15012 N15011 N15012 10
D15012 N15012 0 diode
R15013 N15012 N15013 10
D15013 N15013 0 diode
R15014 N15013 N15014 10
D15014 N15014 0 diode
R15015 N15014 N15015 10
D15015 N15015 0 diode
R15016 N15015 N15016 10
D15016 N15016 0 diode
R15017 N15016 N15017 10
D15017 N15017 0 diode
R15018 N15017 N15018 10
D15018 N15018 0 diode
R15019 N15018 N15019 10
D15019 N15019 0 diode
R15020 N15019 N15020 10
D15020 N15020 0 diode
R15021 N15020 N15021 10
D15021 N15021 0 diode
R15022 N15021 N15022 10
D15022 N15022 0 diode
R15023 N15022 N15023 10
D15023 N15023 0 diode
R15024 N15023 N15024 10
D15024 N15024 0 diode
R15025 N15024 N15025 10
D15025 N15025 0 diode
R15026 N15025 N15026 10
D15026 N15026 0 diode
R15027 N15026 N15027 10
D15027 N15027 0 diode
R15028 N15027 N15028 10
D15028 N15028 0 diode
R15029 N15028 N15029 10
D15029 N15029 0 diode
R15030 N15029 N15030 10
D15030 N15030 0 diode
R15031 N15030 N15031 10
D15031 N15031 0 diode
R15032 N15031 N15032 10
D15032 N15032 0 diode
R15033 N15032 N15033 10
D15033 N15033 0 diode
R15034 N15033 N15034 10
D15034 N15034 0 diode
R15035 N15034 N15035 10
D15035 N15035 0 diode
R15036 N15035 N15036 10
D15036 N15036 0 diode
R15037 N15036 N15037 10
D15037 N15037 0 diode
R15038 N15037 N15038 10
D15038 N15038 0 diode
R15039 N15038 N15039 10
D15039 N15039 0 diode
R15040 N15039 N15040 10
D15040 N15040 0 diode
R15041 N15040 N15041 10
D15041 N15041 0 diode
R15042 N15041 N15042 10
D15042 N15042 0 diode
R15043 N15042 N15043 10
D15043 N15043 0 diode
R15044 N15043 N15044 10
D15044 N15044 0 diode
R15045 N15044 N15045 10
D15045 N15045 0 diode
R15046 N15045 N15046 10
D15046 N15046 0 diode
R15047 N15046 N15047 10
D15047 N15047 0 diode
R15048 N15047 N15048 10
D15048 N15048 0 diode
R15049 N15048 N15049 10
D15049 N15049 0 diode
R15050 N15049 N15050 10
D15050 N15050 0 diode
R15051 N15050 N15051 10
D15051 N15051 0 diode
R15052 N15051 N15052 10
D15052 N15052 0 diode
R15053 N15052 N15053 10
D15053 N15053 0 diode
R15054 N15053 N15054 10
D15054 N15054 0 diode
R15055 N15054 N15055 10
D15055 N15055 0 diode
R15056 N15055 N15056 10
D15056 N15056 0 diode
R15057 N15056 N15057 10
D15057 N15057 0 diode
R15058 N15057 N15058 10
D15058 N15058 0 diode
R15059 N15058 N15059 10
D15059 N15059 0 diode
R15060 N15059 N15060 10
D15060 N15060 0 diode
R15061 N15060 N15061 10
D15061 N15061 0 diode
R15062 N15061 N15062 10
D15062 N15062 0 diode
R15063 N15062 N15063 10
D15063 N15063 0 diode
R15064 N15063 N15064 10
D15064 N15064 0 diode
R15065 N15064 N15065 10
D15065 N15065 0 diode
R15066 N15065 N15066 10
D15066 N15066 0 diode
R15067 N15066 N15067 10
D15067 N15067 0 diode
R15068 N15067 N15068 10
D15068 N15068 0 diode
R15069 N15068 N15069 10
D15069 N15069 0 diode
R15070 N15069 N15070 10
D15070 N15070 0 diode
R15071 N15070 N15071 10
D15071 N15071 0 diode
R15072 N15071 N15072 10
D15072 N15072 0 diode
R15073 N15072 N15073 10
D15073 N15073 0 diode
R15074 N15073 N15074 10
D15074 N15074 0 diode
R15075 N15074 N15075 10
D15075 N15075 0 diode
R15076 N15075 N15076 10
D15076 N15076 0 diode
R15077 N15076 N15077 10
D15077 N15077 0 diode
R15078 N15077 N15078 10
D15078 N15078 0 diode
R15079 N15078 N15079 10
D15079 N15079 0 diode
R15080 N15079 N15080 10
D15080 N15080 0 diode
R15081 N15080 N15081 10
D15081 N15081 0 diode
R15082 N15081 N15082 10
D15082 N15082 0 diode
R15083 N15082 N15083 10
D15083 N15083 0 diode
R15084 N15083 N15084 10
D15084 N15084 0 diode
R15085 N15084 N15085 10
D15085 N15085 0 diode
R15086 N15085 N15086 10
D15086 N15086 0 diode
R15087 N15086 N15087 10
D15087 N15087 0 diode
R15088 N15087 N15088 10
D15088 N15088 0 diode
R15089 N15088 N15089 10
D15089 N15089 0 diode
R15090 N15089 N15090 10
D15090 N15090 0 diode
R15091 N15090 N15091 10
D15091 N15091 0 diode
R15092 N15091 N15092 10
D15092 N15092 0 diode
R15093 N15092 N15093 10
D15093 N15093 0 diode
R15094 N15093 N15094 10
D15094 N15094 0 diode
R15095 N15094 N15095 10
D15095 N15095 0 diode
R15096 N15095 N15096 10
D15096 N15096 0 diode
R15097 N15096 N15097 10
D15097 N15097 0 diode
R15098 N15097 N15098 10
D15098 N15098 0 diode
R15099 N15098 N15099 10
D15099 N15099 0 diode
R15100 N15099 N15100 10
D15100 N15100 0 diode
R15101 N15100 N15101 10
D15101 N15101 0 diode
R15102 N15101 N15102 10
D15102 N15102 0 diode
R15103 N15102 N15103 10
D15103 N15103 0 diode
R15104 N15103 N15104 10
D15104 N15104 0 diode
R15105 N15104 N15105 10
D15105 N15105 0 diode
R15106 N15105 N15106 10
D15106 N15106 0 diode
R15107 N15106 N15107 10
D15107 N15107 0 diode
R15108 N15107 N15108 10
D15108 N15108 0 diode
R15109 N15108 N15109 10
D15109 N15109 0 diode
R15110 N15109 N15110 10
D15110 N15110 0 diode
R15111 N15110 N15111 10
D15111 N15111 0 diode
R15112 N15111 N15112 10
D15112 N15112 0 diode
R15113 N15112 N15113 10
D15113 N15113 0 diode
R15114 N15113 N15114 10
D15114 N15114 0 diode
R15115 N15114 N15115 10
D15115 N15115 0 diode
R15116 N15115 N15116 10
D15116 N15116 0 diode
R15117 N15116 N15117 10
D15117 N15117 0 diode
R15118 N15117 N15118 10
D15118 N15118 0 diode
R15119 N15118 N15119 10
D15119 N15119 0 diode
R15120 N15119 N15120 10
D15120 N15120 0 diode
R15121 N15120 N15121 10
D15121 N15121 0 diode
R15122 N15121 N15122 10
D15122 N15122 0 diode
R15123 N15122 N15123 10
D15123 N15123 0 diode
R15124 N15123 N15124 10
D15124 N15124 0 diode
R15125 N15124 N15125 10
D15125 N15125 0 diode
R15126 N15125 N15126 10
D15126 N15126 0 diode
R15127 N15126 N15127 10
D15127 N15127 0 diode
R15128 N15127 N15128 10
D15128 N15128 0 diode
R15129 N15128 N15129 10
D15129 N15129 0 diode
R15130 N15129 N15130 10
D15130 N15130 0 diode
R15131 N15130 N15131 10
D15131 N15131 0 diode
R15132 N15131 N15132 10
D15132 N15132 0 diode
R15133 N15132 N15133 10
D15133 N15133 0 diode
R15134 N15133 N15134 10
D15134 N15134 0 diode
R15135 N15134 N15135 10
D15135 N15135 0 diode
R15136 N15135 N15136 10
D15136 N15136 0 diode
R15137 N15136 N15137 10
D15137 N15137 0 diode
R15138 N15137 N15138 10
D15138 N15138 0 diode
R15139 N15138 N15139 10
D15139 N15139 0 diode
R15140 N15139 N15140 10
D15140 N15140 0 diode
R15141 N15140 N15141 10
D15141 N15141 0 diode
R15142 N15141 N15142 10
D15142 N15142 0 diode
R15143 N15142 N15143 10
D15143 N15143 0 diode
R15144 N15143 N15144 10
D15144 N15144 0 diode
R15145 N15144 N15145 10
D15145 N15145 0 diode
R15146 N15145 N15146 10
D15146 N15146 0 diode
R15147 N15146 N15147 10
D15147 N15147 0 diode
R15148 N15147 N15148 10
D15148 N15148 0 diode
R15149 N15148 N15149 10
D15149 N15149 0 diode
R15150 N15149 N15150 10
D15150 N15150 0 diode
R15151 N15150 N15151 10
D15151 N15151 0 diode
R15152 N15151 N15152 10
D15152 N15152 0 diode
R15153 N15152 N15153 10
D15153 N15153 0 diode
R15154 N15153 N15154 10
D15154 N15154 0 diode
R15155 N15154 N15155 10
D15155 N15155 0 diode
R15156 N15155 N15156 10
D15156 N15156 0 diode
R15157 N15156 N15157 10
D15157 N15157 0 diode
R15158 N15157 N15158 10
D15158 N15158 0 diode
R15159 N15158 N15159 10
D15159 N15159 0 diode
R15160 N15159 N15160 10
D15160 N15160 0 diode
R15161 N15160 N15161 10
D15161 N15161 0 diode
R15162 N15161 N15162 10
D15162 N15162 0 diode
R15163 N15162 N15163 10
D15163 N15163 0 diode
R15164 N15163 N15164 10
D15164 N15164 0 diode
R15165 N15164 N15165 10
D15165 N15165 0 diode
R15166 N15165 N15166 10
D15166 N15166 0 diode
R15167 N15166 N15167 10
D15167 N15167 0 diode
R15168 N15167 N15168 10
D15168 N15168 0 diode
R15169 N15168 N15169 10
D15169 N15169 0 diode
R15170 N15169 N15170 10
D15170 N15170 0 diode
R15171 N15170 N15171 10
D15171 N15171 0 diode
R15172 N15171 N15172 10
D15172 N15172 0 diode
R15173 N15172 N15173 10
D15173 N15173 0 diode
R15174 N15173 N15174 10
D15174 N15174 0 diode
R15175 N15174 N15175 10
D15175 N15175 0 diode
R15176 N15175 N15176 10
D15176 N15176 0 diode
R15177 N15176 N15177 10
D15177 N15177 0 diode
R15178 N15177 N15178 10
D15178 N15178 0 diode
R15179 N15178 N15179 10
D15179 N15179 0 diode
R15180 N15179 N15180 10
D15180 N15180 0 diode
R15181 N15180 N15181 10
D15181 N15181 0 diode
R15182 N15181 N15182 10
D15182 N15182 0 diode
R15183 N15182 N15183 10
D15183 N15183 0 diode
R15184 N15183 N15184 10
D15184 N15184 0 diode
R15185 N15184 N15185 10
D15185 N15185 0 diode
R15186 N15185 N15186 10
D15186 N15186 0 diode
R15187 N15186 N15187 10
D15187 N15187 0 diode
R15188 N15187 N15188 10
D15188 N15188 0 diode
R15189 N15188 N15189 10
D15189 N15189 0 diode
R15190 N15189 N15190 10
D15190 N15190 0 diode
R15191 N15190 N15191 10
D15191 N15191 0 diode
R15192 N15191 N15192 10
D15192 N15192 0 diode
R15193 N15192 N15193 10
D15193 N15193 0 diode
R15194 N15193 N15194 10
D15194 N15194 0 diode
R15195 N15194 N15195 10
D15195 N15195 0 diode
R15196 N15195 N15196 10
D15196 N15196 0 diode
R15197 N15196 N15197 10
D15197 N15197 0 diode
R15198 N15197 N15198 10
D15198 N15198 0 diode
R15199 N15198 N15199 10
D15199 N15199 0 diode
R15200 N15199 N15200 10
D15200 N15200 0 diode
R15201 N15200 N15201 10
D15201 N15201 0 diode
R15202 N15201 N15202 10
D15202 N15202 0 diode
R15203 N15202 N15203 10
D15203 N15203 0 diode
R15204 N15203 N15204 10
D15204 N15204 0 diode
R15205 N15204 N15205 10
D15205 N15205 0 diode
R15206 N15205 N15206 10
D15206 N15206 0 diode
R15207 N15206 N15207 10
D15207 N15207 0 diode
R15208 N15207 N15208 10
D15208 N15208 0 diode
R15209 N15208 N15209 10
D15209 N15209 0 diode
R15210 N15209 N15210 10
D15210 N15210 0 diode
R15211 N15210 N15211 10
D15211 N15211 0 diode
R15212 N15211 N15212 10
D15212 N15212 0 diode
R15213 N15212 N15213 10
D15213 N15213 0 diode
R15214 N15213 N15214 10
D15214 N15214 0 diode
R15215 N15214 N15215 10
D15215 N15215 0 diode
R15216 N15215 N15216 10
D15216 N15216 0 diode
R15217 N15216 N15217 10
D15217 N15217 0 diode
R15218 N15217 N15218 10
D15218 N15218 0 diode
R15219 N15218 N15219 10
D15219 N15219 0 diode
R15220 N15219 N15220 10
D15220 N15220 0 diode
R15221 N15220 N15221 10
D15221 N15221 0 diode
R15222 N15221 N15222 10
D15222 N15222 0 diode
R15223 N15222 N15223 10
D15223 N15223 0 diode
R15224 N15223 N15224 10
D15224 N15224 0 diode
R15225 N15224 N15225 10
D15225 N15225 0 diode
R15226 N15225 N15226 10
D15226 N15226 0 diode
R15227 N15226 N15227 10
D15227 N15227 0 diode
R15228 N15227 N15228 10
D15228 N15228 0 diode
R15229 N15228 N15229 10
D15229 N15229 0 diode
R15230 N15229 N15230 10
D15230 N15230 0 diode
R15231 N15230 N15231 10
D15231 N15231 0 diode
R15232 N15231 N15232 10
D15232 N15232 0 diode
R15233 N15232 N15233 10
D15233 N15233 0 diode
R15234 N15233 N15234 10
D15234 N15234 0 diode
R15235 N15234 N15235 10
D15235 N15235 0 diode
R15236 N15235 N15236 10
D15236 N15236 0 diode
R15237 N15236 N15237 10
D15237 N15237 0 diode
R15238 N15237 N15238 10
D15238 N15238 0 diode
R15239 N15238 N15239 10
D15239 N15239 0 diode
R15240 N15239 N15240 10
D15240 N15240 0 diode
R15241 N15240 N15241 10
D15241 N15241 0 diode
R15242 N15241 N15242 10
D15242 N15242 0 diode
R15243 N15242 N15243 10
D15243 N15243 0 diode
R15244 N15243 N15244 10
D15244 N15244 0 diode
R15245 N15244 N15245 10
D15245 N15245 0 diode
R15246 N15245 N15246 10
D15246 N15246 0 diode
R15247 N15246 N15247 10
D15247 N15247 0 diode
R15248 N15247 N15248 10
D15248 N15248 0 diode
R15249 N15248 N15249 10
D15249 N15249 0 diode
R15250 N15249 N15250 10
D15250 N15250 0 diode
R15251 N15250 N15251 10
D15251 N15251 0 diode
R15252 N15251 N15252 10
D15252 N15252 0 diode
R15253 N15252 N15253 10
D15253 N15253 0 diode
R15254 N15253 N15254 10
D15254 N15254 0 diode
R15255 N15254 N15255 10
D15255 N15255 0 diode
R15256 N15255 N15256 10
D15256 N15256 0 diode
R15257 N15256 N15257 10
D15257 N15257 0 diode
R15258 N15257 N15258 10
D15258 N15258 0 diode
R15259 N15258 N15259 10
D15259 N15259 0 diode
R15260 N15259 N15260 10
D15260 N15260 0 diode
R15261 N15260 N15261 10
D15261 N15261 0 diode
R15262 N15261 N15262 10
D15262 N15262 0 diode
R15263 N15262 N15263 10
D15263 N15263 0 diode
R15264 N15263 N15264 10
D15264 N15264 0 diode
R15265 N15264 N15265 10
D15265 N15265 0 diode
R15266 N15265 N15266 10
D15266 N15266 0 diode
R15267 N15266 N15267 10
D15267 N15267 0 diode
R15268 N15267 N15268 10
D15268 N15268 0 diode
R15269 N15268 N15269 10
D15269 N15269 0 diode
R15270 N15269 N15270 10
D15270 N15270 0 diode
R15271 N15270 N15271 10
D15271 N15271 0 diode
R15272 N15271 N15272 10
D15272 N15272 0 diode
R15273 N15272 N15273 10
D15273 N15273 0 diode
R15274 N15273 N15274 10
D15274 N15274 0 diode
R15275 N15274 N15275 10
D15275 N15275 0 diode
R15276 N15275 N15276 10
D15276 N15276 0 diode
R15277 N15276 N15277 10
D15277 N15277 0 diode
R15278 N15277 N15278 10
D15278 N15278 0 diode
R15279 N15278 N15279 10
D15279 N15279 0 diode
R15280 N15279 N15280 10
D15280 N15280 0 diode
R15281 N15280 N15281 10
D15281 N15281 0 diode
R15282 N15281 N15282 10
D15282 N15282 0 diode
R15283 N15282 N15283 10
D15283 N15283 0 diode
R15284 N15283 N15284 10
D15284 N15284 0 diode
R15285 N15284 N15285 10
D15285 N15285 0 diode
R15286 N15285 N15286 10
D15286 N15286 0 diode
R15287 N15286 N15287 10
D15287 N15287 0 diode
R15288 N15287 N15288 10
D15288 N15288 0 diode
R15289 N15288 N15289 10
D15289 N15289 0 diode
R15290 N15289 N15290 10
D15290 N15290 0 diode
R15291 N15290 N15291 10
D15291 N15291 0 diode
R15292 N15291 N15292 10
D15292 N15292 0 diode
R15293 N15292 N15293 10
D15293 N15293 0 diode
R15294 N15293 N15294 10
D15294 N15294 0 diode
R15295 N15294 N15295 10
D15295 N15295 0 diode
R15296 N15295 N15296 10
D15296 N15296 0 diode
R15297 N15296 N15297 10
D15297 N15297 0 diode
R15298 N15297 N15298 10
D15298 N15298 0 diode
R15299 N15298 N15299 10
D15299 N15299 0 diode
R15300 N15299 N15300 10
D15300 N15300 0 diode
R15301 N15300 N15301 10
D15301 N15301 0 diode
R15302 N15301 N15302 10
D15302 N15302 0 diode
R15303 N15302 N15303 10
D15303 N15303 0 diode
R15304 N15303 N15304 10
D15304 N15304 0 diode
R15305 N15304 N15305 10
D15305 N15305 0 diode
R15306 N15305 N15306 10
D15306 N15306 0 diode
R15307 N15306 N15307 10
D15307 N15307 0 diode
R15308 N15307 N15308 10
D15308 N15308 0 diode
R15309 N15308 N15309 10
D15309 N15309 0 diode
R15310 N15309 N15310 10
D15310 N15310 0 diode
R15311 N15310 N15311 10
D15311 N15311 0 diode
R15312 N15311 N15312 10
D15312 N15312 0 diode
R15313 N15312 N15313 10
D15313 N15313 0 diode
R15314 N15313 N15314 10
D15314 N15314 0 diode
R15315 N15314 N15315 10
D15315 N15315 0 diode
R15316 N15315 N15316 10
D15316 N15316 0 diode
R15317 N15316 N15317 10
D15317 N15317 0 diode
R15318 N15317 N15318 10
D15318 N15318 0 diode
R15319 N15318 N15319 10
D15319 N15319 0 diode
R15320 N15319 N15320 10
D15320 N15320 0 diode
R15321 N15320 N15321 10
D15321 N15321 0 diode
R15322 N15321 N15322 10
D15322 N15322 0 diode
R15323 N15322 N15323 10
D15323 N15323 0 diode
R15324 N15323 N15324 10
D15324 N15324 0 diode
R15325 N15324 N15325 10
D15325 N15325 0 diode
R15326 N15325 N15326 10
D15326 N15326 0 diode
R15327 N15326 N15327 10
D15327 N15327 0 diode
R15328 N15327 N15328 10
D15328 N15328 0 diode
R15329 N15328 N15329 10
D15329 N15329 0 diode
R15330 N15329 N15330 10
D15330 N15330 0 diode
R15331 N15330 N15331 10
D15331 N15331 0 diode
R15332 N15331 N15332 10
D15332 N15332 0 diode
R15333 N15332 N15333 10
D15333 N15333 0 diode
R15334 N15333 N15334 10
D15334 N15334 0 diode
R15335 N15334 N15335 10
D15335 N15335 0 diode
R15336 N15335 N15336 10
D15336 N15336 0 diode
R15337 N15336 N15337 10
D15337 N15337 0 diode
R15338 N15337 N15338 10
D15338 N15338 0 diode
R15339 N15338 N15339 10
D15339 N15339 0 diode
R15340 N15339 N15340 10
D15340 N15340 0 diode
R15341 N15340 N15341 10
D15341 N15341 0 diode
R15342 N15341 N15342 10
D15342 N15342 0 diode
R15343 N15342 N15343 10
D15343 N15343 0 diode
R15344 N15343 N15344 10
D15344 N15344 0 diode
R15345 N15344 N15345 10
D15345 N15345 0 diode
R15346 N15345 N15346 10
D15346 N15346 0 diode
R15347 N15346 N15347 10
D15347 N15347 0 diode
R15348 N15347 N15348 10
D15348 N15348 0 diode
R15349 N15348 N15349 10
D15349 N15349 0 diode
R15350 N15349 N15350 10
D15350 N15350 0 diode
R15351 N15350 N15351 10
D15351 N15351 0 diode
R15352 N15351 N15352 10
D15352 N15352 0 diode
R15353 N15352 N15353 10
D15353 N15353 0 diode
R15354 N15353 N15354 10
D15354 N15354 0 diode
R15355 N15354 N15355 10
D15355 N15355 0 diode
R15356 N15355 N15356 10
D15356 N15356 0 diode
R15357 N15356 N15357 10
D15357 N15357 0 diode
R15358 N15357 N15358 10
D15358 N15358 0 diode
R15359 N15358 N15359 10
D15359 N15359 0 diode
R15360 N15359 N15360 10
D15360 N15360 0 diode
R15361 N15360 N15361 10
D15361 N15361 0 diode
R15362 N15361 N15362 10
D15362 N15362 0 diode
R15363 N15362 N15363 10
D15363 N15363 0 diode
R15364 N15363 N15364 10
D15364 N15364 0 diode
R15365 N15364 N15365 10
D15365 N15365 0 diode
R15366 N15365 N15366 10
D15366 N15366 0 diode
R15367 N15366 N15367 10
D15367 N15367 0 diode
R15368 N15367 N15368 10
D15368 N15368 0 diode
R15369 N15368 N15369 10
D15369 N15369 0 diode
R15370 N15369 N15370 10
D15370 N15370 0 diode
R15371 N15370 N15371 10
D15371 N15371 0 diode
R15372 N15371 N15372 10
D15372 N15372 0 diode
R15373 N15372 N15373 10
D15373 N15373 0 diode
R15374 N15373 N15374 10
D15374 N15374 0 diode
R15375 N15374 N15375 10
D15375 N15375 0 diode
R15376 N15375 N15376 10
D15376 N15376 0 diode
R15377 N15376 N15377 10
D15377 N15377 0 diode
R15378 N15377 N15378 10
D15378 N15378 0 diode
R15379 N15378 N15379 10
D15379 N15379 0 diode
R15380 N15379 N15380 10
D15380 N15380 0 diode
R15381 N15380 N15381 10
D15381 N15381 0 diode
R15382 N15381 N15382 10
D15382 N15382 0 diode
R15383 N15382 N15383 10
D15383 N15383 0 diode
R15384 N15383 N15384 10
D15384 N15384 0 diode
R15385 N15384 N15385 10
D15385 N15385 0 diode
R15386 N15385 N15386 10
D15386 N15386 0 diode
R15387 N15386 N15387 10
D15387 N15387 0 diode
R15388 N15387 N15388 10
D15388 N15388 0 diode
R15389 N15388 N15389 10
D15389 N15389 0 diode
R15390 N15389 N15390 10
D15390 N15390 0 diode
R15391 N15390 N15391 10
D15391 N15391 0 diode
R15392 N15391 N15392 10
D15392 N15392 0 diode
R15393 N15392 N15393 10
D15393 N15393 0 diode
R15394 N15393 N15394 10
D15394 N15394 0 diode
R15395 N15394 N15395 10
D15395 N15395 0 diode
R15396 N15395 N15396 10
D15396 N15396 0 diode
R15397 N15396 N15397 10
D15397 N15397 0 diode
R15398 N15397 N15398 10
D15398 N15398 0 diode
R15399 N15398 N15399 10
D15399 N15399 0 diode
R15400 N15399 N15400 10
D15400 N15400 0 diode
R15401 N15400 N15401 10
D15401 N15401 0 diode
R15402 N15401 N15402 10
D15402 N15402 0 diode
R15403 N15402 N15403 10
D15403 N15403 0 diode
R15404 N15403 N15404 10
D15404 N15404 0 diode
R15405 N15404 N15405 10
D15405 N15405 0 diode
R15406 N15405 N15406 10
D15406 N15406 0 diode
R15407 N15406 N15407 10
D15407 N15407 0 diode
R15408 N15407 N15408 10
D15408 N15408 0 diode
R15409 N15408 N15409 10
D15409 N15409 0 diode
R15410 N15409 N15410 10
D15410 N15410 0 diode
R15411 N15410 N15411 10
D15411 N15411 0 diode
R15412 N15411 N15412 10
D15412 N15412 0 diode
R15413 N15412 N15413 10
D15413 N15413 0 diode
R15414 N15413 N15414 10
D15414 N15414 0 diode
R15415 N15414 N15415 10
D15415 N15415 0 diode
R15416 N15415 N15416 10
D15416 N15416 0 diode
R15417 N15416 N15417 10
D15417 N15417 0 diode
R15418 N15417 N15418 10
D15418 N15418 0 diode
R15419 N15418 N15419 10
D15419 N15419 0 diode
R15420 N15419 N15420 10
D15420 N15420 0 diode
R15421 N15420 N15421 10
D15421 N15421 0 diode
R15422 N15421 N15422 10
D15422 N15422 0 diode
R15423 N15422 N15423 10
D15423 N15423 0 diode
R15424 N15423 N15424 10
D15424 N15424 0 diode
R15425 N15424 N15425 10
D15425 N15425 0 diode
R15426 N15425 N15426 10
D15426 N15426 0 diode
R15427 N15426 N15427 10
D15427 N15427 0 diode
R15428 N15427 N15428 10
D15428 N15428 0 diode
R15429 N15428 N15429 10
D15429 N15429 0 diode
R15430 N15429 N15430 10
D15430 N15430 0 diode
R15431 N15430 N15431 10
D15431 N15431 0 diode
R15432 N15431 N15432 10
D15432 N15432 0 diode
R15433 N15432 N15433 10
D15433 N15433 0 diode
R15434 N15433 N15434 10
D15434 N15434 0 diode
R15435 N15434 N15435 10
D15435 N15435 0 diode
R15436 N15435 N15436 10
D15436 N15436 0 diode
R15437 N15436 N15437 10
D15437 N15437 0 diode
R15438 N15437 N15438 10
D15438 N15438 0 diode
R15439 N15438 N15439 10
D15439 N15439 0 diode
R15440 N15439 N15440 10
D15440 N15440 0 diode
R15441 N15440 N15441 10
D15441 N15441 0 diode
R15442 N15441 N15442 10
D15442 N15442 0 diode
R15443 N15442 N15443 10
D15443 N15443 0 diode
R15444 N15443 N15444 10
D15444 N15444 0 diode
R15445 N15444 N15445 10
D15445 N15445 0 diode
R15446 N15445 N15446 10
D15446 N15446 0 diode
R15447 N15446 N15447 10
D15447 N15447 0 diode
R15448 N15447 N15448 10
D15448 N15448 0 diode
R15449 N15448 N15449 10
D15449 N15449 0 diode
R15450 N15449 N15450 10
D15450 N15450 0 diode
R15451 N15450 N15451 10
D15451 N15451 0 diode
R15452 N15451 N15452 10
D15452 N15452 0 diode
R15453 N15452 N15453 10
D15453 N15453 0 diode
R15454 N15453 N15454 10
D15454 N15454 0 diode
R15455 N15454 N15455 10
D15455 N15455 0 diode
R15456 N15455 N15456 10
D15456 N15456 0 diode
R15457 N15456 N15457 10
D15457 N15457 0 diode
R15458 N15457 N15458 10
D15458 N15458 0 diode
R15459 N15458 N15459 10
D15459 N15459 0 diode
R15460 N15459 N15460 10
D15460 N15460 0 diode
R15461 N15460 N15461 10
D15461 N15461 0 diode
R15462 N15461 N15462 10
D15462 N15462 0 diode
R15463 N15462 N15463 10
D15463 N15463 0 diode
R15464 N15463 N15464 10
D15464 N15464 0 diode
R15465 N15464 N15465 10
D15465 N15465 0 diode
R15466 N15465 N15466 10
D15466 N15466 0 diode
R15467 N15466 N15467 10
D15467 N15467 0 diode
R15468 N15467 N15468 10
D15468 N15468 0 diode
R15469 N15468 N15469 10
D15469 N15469 0 diode
R15470 N15469 N15470 10
D15470 N15470 0 diode
R15471 N15470 N15471 10
D15471 N15471 0 diode
R15472 N15471 N15472 10
D15472 N15472 0 diode
R15473 N15472 N15473 10
D15473 N15473 0 diode
R15474 N15473 N15474 10
D15474 N15474 0 diode
R15475 N15474 N15475 10
D15475 N15475 0 diode
R15476 N15475 N15476 10
D15476 N15476 0 diode
R15477 N15476 N15477 10
D15477 N15477 0 diode
R15478 N15477 N15478 10
D15478 N15478 0 diode
R15479 N15478 N15479 10
D15479 N15479 0 diode
R15480 N15479 N15480 10
D15480 N15480 0 diode
R15481 N15480 N15481 10
D15481 N15481 0 diode
R15482 N15481 N15482 10
D15482 N15482 0 diode
R15483 N15482 N15483 10
D15483 N15483 0 diode
R15484 N15483 N15484 10
D15484 N15484 0 diode
R15485 N15484 N15485 10
D15485 N15485 0 diode
R15486 N15485 N15486 10
D15486 N15486 0 diode
R15487 N15486 N15487 10
D15487 N15487 0 diode
R15488 N15487 N15488 10
D15488 N15488 0 diode
R15489 N15488 N15489 10
D15489 N15489 0 diode
R15490 N15489 N15490 10
D15490 N15490 0 diode
R15491 N15490 N15491 10
D15491 N15491 0 diode
R15492 N15491 N15492 10
D15492 N15492 0 diode
R15493 N15492 N15493 10
D15493 N15493 0 diode
R15494 N15493 N15494 10
D15494 N15494 0 diode
R15495 N15494 N15495 10
D15495 N15495 0 diode
R15496 N15495 N15496 10
D15496 N15496 0 diode
R15497 N15496 N15497 10
D15497 N15497 0 diode
R15498 N15497 N15498 10
D15498 N15498 0 diode
R15499 N15498 N15499 10
D15499 N15499 0 diode
R15500 N15499 N15500 10
D15500 N15500 0 diode
R15501 N15500 N15501 10
D15501 N15501 0 diode
R15502 N15501 N15502 10
D15502 N15502 0 diode
R15503 N15502 N15503 10
D15503 N15503 0 diode
R15504 N15503 N15504 10
D15504 N15504 0 diode
R15505 N15504 N15505 10
D15505 N15505 0 diode
R15506 N15505 N15506 10
D15506 N15506 0 diode
R15507 N15506 N15507 10
D15507 N15507 0 diode
R15508 N15507 N15508 10
D15508 N15508 0 diode
R15509 N15508 N15509 10
D15509 N15509 0 diode
R15510 N15509 N15510 10
D15510 N15510 0 diode
R15511 N15510 N15511 10
D15511 N15511 0 diode
R15512 N15511 N15512 10
D15512 N15512 0 diode
R15513 N15512 N15513 10
D15513 N15513 0 diode
R15514 N15513 N15514 10
D15514 N15514 0 diode
R15515 N15514 N15515 10
D15515 N15515 0 diode
R15516 N15515 N15516 10
D15516 N15516 0 diode
R15517 N15516 N15517 10
D15517 N15517 0 diode
R15518 N15517 N15518 10
D15518 N15518 0 diode
R15519 N15518 N15519 10
D15519 N15519 0 diode
R15520 N15519 N15520 10
D15520 N15520 0 diode
R15521 N15520 N15521 10
D15521 N15521 0 diode
R15522 N15521 N15522 10
D15522 N15522 0 diode
R15523 N15522 N15523 10
D15523 N15523 0 diode
R15524 N15523 N15524 10
D15524 N15524 0 diode
R15525 N15524 N15525 10
D15525 N15525 0 diode
R15526 N15525 N15526 10
D15526 N15526 0 diode
R15527 N15526 N15527 10
D15527 N15527 0 diode
R15528 N15527 N15528 10
D15528 N15528 0 diode
R15529 N15528 N15529 10
D15529 N15529 0 diode
R15530 N15529 N15530 10
D15530 N15530 0 diode
R15531 N15530 N15531 10
D15531 N15531 0 diode
R15532 N15531 N15532 10
D15532 N15532 0 diode
R15533 N15532 N15533 10
D15533 N15533 0 diode
R15534 N15533 N15534 10
D15534 N15534 0 diode
R15535 N15534 N15535 10
D15535 N15535 0 diode
R15536 N15535 N15536 10
D15536 N15536 0 diode
R15537 N15536 N15537 10
D15537 N15537 0 diode
R15538 N15537 N15538 10
D15538 N15538 0 diode
R15539 N15538 N15539 10
D15539 N15539 0 diode
R15540 N15539 N15540 10
D15540 N15540 0 diode
R15541 N15540 N15541 10
D15541 N15541 0 diode
R15542 N15541 N15542 10
D15542 N15542 0 diode
R15543 N15542 N15543 10
D15543 N15543 0 diode
R15544 N15543 N15544 10
D15544 N15544 0 diode
R15545 N15544 N15545 10
D15545 N15545 0 diode
R15546 N15545 N15546 10
D15546 N15546 0 diode
R15547 N15546 N15547 10
D15547 N15547 0 diode
R15548 N15547 N15548 10
D15548 N15548 0 diode
R15549 N15548 N15549 10
D15549 N15549 0 diode
R15550 N15549 N15550 10
D15550 N15550 0 diode
R15551 N15550 N15551 10
D15551 N15551 0 diode
R15552 N15551 N15552 10
D15552 N15552 0 diode
R15553 N15552 N15553 10
D15553 N15553 0 diode
R15554 N15553 N15554 10
D15554 N15554 0 diode
R15555 N15554 N15555 10
D15555 N15555 0 diode
R15556 N15555 N15556 10
D15556 N15556 0 diode
R15557 N15556 N15557 10
D15557 N15557 0 diode
R15558 N15557 N15558 10
D15558 N15558 0 diode
R15559 N15558 N15559 10
D15559 N15559 0 diode
R15560 N15559 N15560 10
D15560 N15560 0 diode
R15561 N15560 N15561 10
D15561 N15561 0 diode
R15562 N15561 N15562 10
D15562 N15562 0 diode
R15563 N15562 N15563 10
D15563 N15563 0 diode
R15564 N15563 N15564 10
D15564 N15564 0 diode
R15565 N15564 N15565 10
D15565 N15565 0 diode
R15566 N15565 N15566 10
D15566 N15566 0 diode
R15567 N15566 N15567 10
D15567 N15567 0 diode
R15568 N15567 N15568 10
D15568 N15568 0 diode
R15569 N15568 N15569 10
D15569 N15569 0 diode
R15570 N15569 N15570 10
D15570 N15570 0 diode
R15571 N15570 N15571 10
D15571 N15571 0 diode
R15572 N15571 N15572 10
D15572 N15572 0 diode
R15573 N15572 N15573 10
D15573 N15573 0 diode
R15574 N15573 N15574 10
D15574 N15574 0 diode
R15575 N15574 N15575 10
D15575 N15575 0 diode
R15576 N15575 N15576 10
D15576 N15576 0 diode
R15577 N15576 N15577 10
D15577 N15577 0 diode
R15578 N15577 N15578 10
D15578 N15578 0 diode
R15579 N15578 N15579 10
D15579 N15579 0 diode
R15580 N15579 N15580 10
D15580 N15580 0 diode
R15581 N15580 N15581 10
D15581 N15581 0 diode
R15582 N15581 N15582 10
D15582 N15582 0 diode
R15583 N15582 N15583 10
D15583 N15583 0 diode
R15584 N15583 N15584 10
D15584 N15584 0 diode
R15585 N15584 N15585 10
D15585 N15585 0 diode
R15586 N15585 N15586 10
D15586 N15586 0 diode
R15587 N15586 N15587 10
D15587 N15587 0 diode
R15588 N15587 N15588 10
D15588 N15588 0 diode
R15589 N15588 N15589 10
D15589 N15589 0 diode
R15590 N15589 N15590 10
D15590 N15590 0 diode
R15591 N15590 N15591 10
D15591 N15591 0 diode
R15592 N15591 N15592 10
D15592 N15592 0 diode
R15593 N15592 N15593 10
D15593 N15593 0 diode
R15594 N15593 N15594 10
D15594 N15594 0 diode
R15595 N15594 N15595 10
D15595 N15595 0 diode
R15596 N15595 N15596 10
D15596 N15596 0 diode
R15597 N15596 N15597 10
D15597 N15597 0 diode
R15598 N15597 N15598 10
D15598 N15598 0 diode
R15599 N15598 N15599 10
D15599 N15599 0 diode
R15600 N15599 N15600 10
D15600 N15600 0 diode
R15601 N15600 N15601 10
D15601 N15601 0 diode
R15602 N15601 N15602 10
D15602 N15602 0 diode
R15603 N15602 N15603 10
D15603 N15603 0 diode
R15604 N15603 N15604 10
D15604 N15604 0 diode
R15605 N15604 N15605 10
D15605 N15605 0 diode
R15606 N15605 N15606 10
D15606 N15606 0 diode
R15607 N15606 N15607 10
D15607 N15607 0 diode
R15608 N15607 N15608 10
D15608 N15608 0 diode
R15609 N15608 N15609 10
D15609 N15609 0 diode
R15610 N15609 N15610 10
D15610 N15610 0 diode
R15611 N15610 N15611 10
D15611 N15611 0 diode
R15612 N15611 N15612 10
D15612 N15612 0 diode
R15613 N15612 N15613 10
D15613 N15613 0 diode
R15614 N15613 N15614 10
D15614 N15614 0 diode
R15615 N15614 N15615 10
D15615 N15615 0 diode
R15616 N15615 N15616 10
D15616 N15616 0 diode
R15617 N15616 N15617 10
D15617 N15617 0 diode
R15618 N15617 N15618 10
D15618 N15618 0 diode
R15619 N15618 N15619 10
D15619 N15619 0 diode
R15620 N15619 N15620 10
D15620 N15620 0 diode
R15621 N15620 N15621 10
D15621 N15621 0 diode
R15622 N15621 N15622 10
D15622 N15622 0 diode
R15623 N15622 N15623 10
D15623 N15623 0 diode
R15624 N15623 N15624 10
D15624 N15624 0 diode
R15625 N15624 N15625 10
D15625 N15625 0 diode
R15626 N15625 N15626 10
D15626 N15626 0 diode
R15627 N15626 N15627 10
D15627 N15627 0 diode
R15628 N15627 N15628 10
D15628 N15628 0 diode
R15629 N15628 N15629 10
D15629 N15629 0 diode
R15630 N15629 N15630 10
D15630 N15630 0 diode
R15631 N15630 N15631 10
D15631 N15631 0 diode
R15632 N15631 N15632 10
D15632 N15632 0 diode
R15633 N15632 N15633 10
D15633 N15633 0 diode
R15634 N15633 N15634 10
D15634 N15634 0 diode
R15635 N15634 N15635 10
D15635 N15635 0 diode
R15636 N15635 N15636 10
D15636 N15636 0 diode
R15637 N15636 N15637 10
D15637 N15637 0 diode
R15638 N15637 N15638 10
D15638 N15638 0 diode
R15639 N15638 N15639 10
D15639 N15639 0 diode
R15640 N15639 N15640 10
D15640 N15640 0 diode
R15641 N15640 N15641 10
D15641 N15641 0 diode
R15642 N15641 N15642 10
D15642 N15642 0 diode
R15643 N15642 N15643 10
D15643 N15643 0 diode
R15644 N15643 N15644 10
D15644 N15644 0 diode
R15645 N15644 N15645 10
D15645 N15645 0 diode
R15646 N15645 N15646 10
D15646 N15646 0 diode
R15647 N15646 N15647 10
D15647 N15647 0 diode
R15648 N15647 N15648 10
D15648 N15648 0 diode
R15649 N15648 N15649 10
D15649 N15649 0 diode
R15650 N15649 N15650 10
D15650 N15650 0 diode
R15651 N15650 N15651 10
D15651 N15651 0 diode
R15652 N15651 N15652 10
D15652 N15652 0 diode
R15653 N15652 N15653 10
D15653 N15653 0 diode
R15654 N15653 N15654 10
D15654 N15654 0 diode
R15655 N15654 N15655 10
D15655 N15655 0 diode
R15656 N15655 N15656 10
D15656 N15656 0 diode
R15657 N15656 N15657 10
D15657 N15657 0 diode
R15658 N15657 N15658 10
D15658 N15658 0 diode
R15659 N15658 N15659 10
D15659 N15659 0 diode
R15660 N15659 N15660 10
D15660 N15660 0 diode
R15661 N15660 N15661 10
D15661 N15661 0 diode
R15662 N15661 N15662 10
D15662 N15662 0 diode
R15663 N15662 N15663 10
D15663 N15663 0 diode
R15664 N15663 N15664 10
D15664 N15664 0 diode
R15665 N15664 N15665 10
D15665 N15665 0 diode
R15666 N15665 N15666 10
D15666 N15666 0 diode
R15667 N15666 N15667 10
D15667 N15667 0 diode
R15668 N15667 N15668 10
D15668 N15668 0 diode
R15669 N15668 N15669 10
D15669 N15669 0 diode
R15670 N15669 N15670 10
D15670 N15670 0 diode
R15671 N15670 N15671 10
D15671 N15671 0 diode
R15672 N15671 N15672 10
D15672 N15672 0 diode
R15673 N15672 N15673 10
D15673 N15673 0 diode
R15674 N15673 N15674 10
D15674 N15674 0 diode
R15675 N15674 N15675 10
D15675 N15675 0 diode
R15676 N15675 N15676 10
D15676 N15676 0 diode
R15677 N15676 N15677 10
D15677 N15677 0 diode
R15678 N15677 N15678 10
D15678 N15678 0 diode
R15679 N15678 N15679 10
D15679 N15679 0 diode
R15680 N15679 N15680 10
D15680 N15680 0 diode
R15681 N15680 N15681 10
D15681 N15681 0 diode
R15682 N15681 N15682 10
D15682 N15682 0 diode
R15683 N15682 N15683 10
D15683 N15683 0 diode
R15684 N15683 N15684 10
D15684 N15684 0 diode
R15685 N15684 N15685 10
D15685 N15685 0 diode
R15686 N15685 N15686 10
D15686 N15686 0 diode
R15687 N15686 N15687 10
D15687 N15687 0 diode
R15688 N15687 N15688 10
D15688 N15688 0 diode
R15689 N15688 N15689 10
D15689 N15689 0 diode
R15690 N15689 N15690 10
D15690 N15690 0 diode
R15691 N15690 N15691 10
D15691 N15691 0 diode
R15692 N15691 N15692 10
D15692 N15692 0 diode
R15693 N15692 N15693 10
D15693 N15693 0 diode
R15694 N15693 N15694 10
D15694 N15694 0 diode
R15695 N15694 N15695 10
D15695 N15695 0 diode
R15696 N15695 N15696 10
D15696 N15696 0 diode
R15697 N15696 N15697 10
D15697 N15697 0 diode
R15698 N15697 N15698 10
D15698 N15698 0 diode
R15699 N15698 N15699 10
D15699 N15699 0 diode
R15700 N15699 N15700 10
D15700 N15700 0 diode
R15701 N15700 N15701 10
D15701 N15701 0 diode
R15702 N15701 N15702 10
D15702 N15702 0 diode
R15703 N15702 N15703 10
D15703 N15703 0 diode
R15704 N15703 N15704 10
D15704 N15704 0 diode
R15705 N15704 N15705 10
D15705 N15705 0 diode
R15706 N15705 N15706 10
D15706 N15706 0 diode
R15707 N15706 N15707 10
D15707 N15707 0 diode
R15708 N15707 N15708 10
D15708 N15708 0 diode
R15709 N15708 N15709 10
D15709 N15709 0 diode
R15710 N15709 N15710 10
D15710 N15710 0 diode
R15711 N15710 N15711 10
D15711 N15711 0 diode
R15712 N15711 N15712 10
D15712 N15712 0 diode
R15713 N15712 N15713 10
D15713 N15713 0 diode
R15714 N15713 N15714 10
D15714 N15714 0 diode
R15715 N15714 N15715 10
D15715 N15715 0 diode
R15716 N15715 N15716 10
D15716 N15716 0 diode
R15717 N15716 N15717 10
D15717 N15717 0 diode
R15718 N15717 N15718 10
D15718 N15718 0 diode
R15719 N15718 N15719 10
D15719 N15719 0 diode
R15720 N15719 N15720 10
D15720 N15720 0 diode
R15721 N15720 N15721 10
D15721 N15721 0 diode
R15722 N15721 N15722 10
D15722 N15722 0 diode
R15723 N15722 N15723 10
D15723 N15723 0 diode
R15724 N15723 N15724 10
D15724 N15724 0 diode
R15725 N15724 N15725 10
D15725 N15725 0 diode
R15726 N15725 N15726 10
D15726 N15726 0 diode
R15727 N15726 N15727 10
D15727 N15727 0 diode
R15728 N15727 N15728 10
D15728 N15728 0 diode
R15729 N15728 N15729 10
D15729 N15729 0 diode
R15730 N15729 N15730 10
D15730 N15730 0 diode
R15731 N15730 N15731 10
D15731 N15731 0 diode
R15732 N15731 N15732 10
D15732 N15732 0 diode
R15733 N15732 N15733 10
D15733 N15733 0 diode
R15734 N15733 N15734 10
D15734 N15734 0 diode
R15735 N15734 N15735 10
D15735 N15735 0 diode
R15736 N15735 N15736 10
D15736 N15736 0 diode
R15737 N15736 N15737 10
D15737 N15737 0 diode
R15738 N15737 N15738 10
D15738 N15738 0 diode
R15739 N15738 N15739 10
D15739 N15739 0 diode
R15740 N15739 N15740 10
D15740 N15740 0 diode
R15741 N15740 N15741 10
D15741 N15741 0 diode
R15742 N15741 N15742 10
D15742 N15742 0 diode
R15743 N15742 N15743 10
D15743 N15743 0 diode
R15744 N15743 N15744 10
D15744 N15744 0 diode
R15745 N15744 N15745 10
D15745 N15745 0 diode
R15746 N15745 N15746 10
D15746 N15746 0 diode
R15747 N15746 N15747 10
D15747 N15747 0 diode
R15748 N15747 N15748 10
D15748 N15748 0 diode
R15749 N15748 N15749 10
D15749 N15749 0 diode
R15750 N15749 N15750 10
D15750 N15750 0 diode
R15751 N15750 N15751 10
D15751 N15751 0 diode
R15752 N15751 N15752 10
D15752 N15752 0 diode
R15753 N15752 N15753 10
D15753 N15753 0 diode
R15754 N15753 N15754 10
D15754 N15754 0 diode
R15755 N15754 N15755 10
D15755 N15755 0 diode
R15756 N15755 N15756 10
D15756 N15756 0 diode
R15757 N15756 N15757 10
D15757 N15757 0 diode
R15758 N15757 N15758 10
D15758 N15758 0 diode
R15759 N15758 N15759 10
D15759 N15759 0 diode
R15760 N15759 N15760 10
D15760 N15760 0 diode
R15761 N15760 N15761 10
D15761 N15761 0 diode
R15762 N15761 N15762 10
D15762 N15762 0 diode
R15763 N15762 N15763 10
D15763 N15763 0 diode
R15764 N15763 N15764 10
D15764 N15764 0 diode
R15765 N15764 N15765 10
D15765 N15765 0 diode
R15766 N15765 N15766 10
D15766 N15766 0 diode
R15767 N15766 N15767 10
D15767 N15767 0 diode
R15768 N15767 N15768 10
D15768 N15768 0 diode
R15769 N15768 N15769 10
D15769 N15769 0 diode
R15770 N15769 N15770 10
D15770 N15770 0 diode
R15771 N15770 N15771 10
D15771 N15771 0 diode
R15772 N15771 N15772 10
D15772 N15772 0 diode
R15773 N15772 N15773 10
D15773 N15773 0 diode
R15774 N15773 N15774 10
D15774 N15774 0 diode
R15775 N15774 N15775 10
D15775 N15775 0 diode
R15776 N15775 N15776 10
D15776 N15776 0 diode
R15777 N15776 N15777 10
D15777 N15777 0 diode
R15778 N15777 N15778 10
D15778 N15778 0 diode
R15779 N15778 N15779 10
D15779 N15779 0 diode
R15780 N15779 N15780 10
D15780 N15780 0 diode
R15781 N15780 N15781 10
D15781 N15781 0 diode
R15782 N15781 N15782 10
D15782 N15782 0 diode
R15783 N15782 N15783 10
D15783 N15783 0 diode
R15784 N15783 N15784 10
D15784 N15784 0 diode
R15785 N15784 N15785 10
D15785 N15785 0 diode
R15786 N15785 N15786 10
D15786 N15786 0 diode
R15787 N15786 N15787 10
D15787 N15787 0 diode
R15788 N15787 N15788 10
D15788 N15788 0 diode
R15789 N15788 N15789 10
D15789 N15789 0 diode
R15790 N15789 N15790 10
D15790 N15790 0 diode
R15791 N15790 N15791 10
D15791 N15791 0 diode
R15792 N15791 N15792 10
D15792 N15792 0 diode
R15793 N15792 N15793 10
D15793 N15793 0 diode
R15794 N15793 N15794 10
D15794 N15794 0 diode
R15795 N15794 N15795 10
D15795 N15795 0 diode
R15796 N15795 N15796 10
D15796 N15796 0 diode
R15797 N15796 N15797 10
D15797 N15797 0 diode
R15798 N15797 N15798 10
D15798 N15798 0 diode
R15799 N15798 N15799 10
D15799 N15799 0 diode
R15800 N15799 N15800 10
D15800 N15800 0 diode
R15801 N15800 N15801 10
D15801 N15801 0 diode
R15802 N15801 N15802 10
D15802 N15802 0 diode
R15803 N15802 N15803 10
D15803 N15803 0 diode
R15804 N15803 N15804 10
D15804 N15804 0 diode
R15805 N15804 N15805 10
D15805 N15805 0 diode
R15806 N15805 N15806 10
D15806 N15806 0 diode
R15807 N15806 N15807 10
D15807 N15807 0 diode
R15808 N15807 N15808 10
D15808 N15808 0 diode
R15809 N15808 N15809 10
D15809 N15809 0 diode
R15810 N15809 N15810 10
D15810 N15810 0 diode
R15811 N15810 N15811 10
D15811 N15811 0 diode
R15812 N15811 N15812 10
D15812 N15812 0 diode
R15813 N15812 N15813 10
D15813 N15813 0 diode
R15814 N15813 N15814 10
D15814 N15814 0 diode
R15815 N15814 N15815 10
D15815 N15815 0 diode
R15816 N15815 N15816 10
D15816 N15816 0 diode
R15817 N15816 N15817 10
D15817 N15817 0 diode
R15818 N15817 N15818 10
D15818 N15818 0 diode
R15819 N15818 N15819 10
D15819 N15819 0 diode
R15820 N15819 N15820 10
D15820 N15820 0 diode
R15821 N15820 N15821 10
D15821 N15821 0 diode
R15822 N15821 N15822 10
D15822 N15822 0 diode
R15823 N15822 N15823 10
D15823 N15823 0 diode
R15824 N15823 N15824 10
D15824 N15824 0 diode
R15825 N15824 N15825 10
D15825 N15825 0 diode
R15826 N15825 N15826 10
D15826 N15826 0 diode
R15827 N15826 N15827 10
D15827 N15827 0 diode
R15828 N15827 N15828 10
D15828 N15828 0 diode
R15829 N15828 N15829 10
D15829 N15829 0 diode
R15830 N15829 N15830 10
D15830 N15830 0 diode
R15831 N15830 N15831 10
D15831 N15831 0 diode
R15832 N15831 N15832 10
D15832 N15832 0 diode
R15833 N15832 N15833 10
D15833 N15833 0 diode
R15834 N15833 N15834 10
D15834 N15834 0 diode
R15835 N15834 N15835 10
D15835 N15835 0 diode
R15836 N15835 N15836 10
D15836 N15836 0 diode
R15837 N15836 N15837 10
D15837 N15837 0 diode
R15838 N15837 N15838 10
D15838 N15838 0 diode
R15839 N15838 N15839 10
D15839 N15839 0 diode
R15840 N15839 N15840 10
D15840 N15840 0 diode
R15841 N15840 N15841 10
D15841 N15841 0 diode
R15842 N15841 N15842 10
D15842 N15842 0 diode
R15843 N15842 N15843 10
D15843 N15843 0 diode
R15844 N15843 N15844 10
D15844 N15844 0 diode
R15845 N15844 N15845 10
D15845 N15845 0 diode
R15846 N15845 N15846 10
D15846 N15846 0 diode
R15847 N15846 N15847 10
D15847 N15847 0 diode
R15848 N15847 N15848 10
D15848 N15848 0 diode
R15849 N15848 N15849 10
D15849 N15849 0 diode
R15850 N15849 N15850 10
D15850 N15850 0 diode
R15851 N15850 N15851 10
D15851 N15851 0 diode
R15852 N15851 N15852 10
D15852 N15852 0 diode
R15853 N15852 N15853 10
D15853 N15853 0 diode
R15854 N15853 N15854 10
D15854 N15854 0 diode
R15855 N15854 N15855 10
D15855 N15855 0 diode
R15856 N15855 N15856 10
D15856 N15856 0 diode
R15857 N15856 N15857 10
D15857 N15857 0 diode
R15858 N15857 N15858 10
D15858 N15858 0 diode
R15859 N15858 N15859 10
D15859 N15859 0 diode
R15860 N15859 N15860 10
D15860 N15860 0 diode
R15861 N15860 N15861 10
D15861 N15861 0 diode
R15862 N15861 N15862 10
D15862 N15862 0 diode
R15863 N15862 N15863 10
D15863 N15863 0 diode
R15864 N15863 N15864 10
D15864 N15864 0 diode
R15865 N15864 N15865 10
D15865 N15865 0 diode
R15866 N15865 N15866 10
D15866 N15866 0 diode
R15867 N15866 N15867 10
D15867 N15867 0 diode
R15868 N15867 N15868 10
D15868 N15868 0 diode
R15869 N15868 N15869 10
D15869 N15869 0 diode
R15870 N15869 N15870 10
D15870 N15870 0 diode
R15871 N15870 N15871 10
D15871 N15871 0 diode
R15872 N15871 N15872 10
D15872 N15872 0 diode
R15873 N15872 N15873 10
D15873 N15873 0 diode
R15874 N15873 N15874 10
D15874 N15874 0 diode
R15875 N15874 N15875 10
D15875 N15875 0 diode
R15876 N15875 N15876 10
D15876 N15876 0 diode
R15877 N15876 N15877 10
D15877 N15877 0 diode
R15878 N15877 N15878 10
D15878 N15878 0 diode
R15879 N15878 N15879 10
D15879 N15879 0 diode
R15880 N15879 N15880 10
D15880 N15880 0 diode
R15881 N15880 N15881 10
D15881 N15881 0 diode
R15882 N15881 N15882 10
D15882 N15882 0 diode
R15883 N15882 N15883 10
D15883 N15883 0 diode
R15884 N15883 N15884 10
D15884 N15884 0 diode
R15885 N15884 N15885 10
D15885 N15885 0 diode
R15886 N15885 N15886 10
D15886 N15886 0 diode
R15887 N15886 N15887 10
D15887 N15887 0 diode
R15888 N15887 N15888 10
D15888 N15888 0 diode
R15889 N15888 N15889 10
D15889 N15889 0 diode
R15890 N15889 N15890 10
D15890 N15890 0 diode
R15891 N15890 N15891 10
D15891 N15891 0 diode
R15892 N15891 N15892 10
D15892 N15892 0 diode
R15893 N15892 N15893 10
D15893 N15893 0 diode
R15894 N15893 N15894 10
D15894 N15894 0 diode
R15895 N15894 N15895 10
D15895 N15895 0 diode
R15896 N15895 N15896 10
D15896 N15896 0 diode
R15897 N15896 N15897 10
D15897 N15897 0 diode
R15898 N15897 N15898 10
D15898 N15898 0 diode
R15899 N15898 N15899 10
D15899 N15899 0 diode
R15900 N15899 N15900 10
D15900 N15900 0 diode
R15901 N15900 N15901 10
D15901 N15901 0 diode
R15902 N15901 N15902 10
D15902 N15902 0 diode
R15903 N15902 N15903 10
D15903 N15903 0 diode
R15904 N15903 N15904 10
D15904 N15904 0 diode
R15905 N15904 N15905 10
D15905 N15905 0 diode
R15906 N15905 N15906 10
D15906 N15906 0 diode
R15907 N15906 N15907 10
D15907 N15907 0 diode
R15908 N15907 N15908 10
D15908 N15908 0 diode
R15909 N15908 N15909 10
D15909 N15909 0 diode
R15910 N15909 N15910 10
D15910 N15910 0 diode
R15911 N15910 N15911 10
D15911 N15911 0 diode
R15912 N15911 N15912 10
D15912 N15912 0 diode
R15913 N15912 N15913 10
D15913 N15913 0 diode
R15914 N15913 N15914 10
D15914 N15914 0 diode
R15915 N15914 N15915 10
D15915 N15915 0 diode
R15916 N15915 N15916 10
D15916 N15916 0 diode
R15917 N15916 N15917 10
D15917 N15917 0 diode
R15918 N15917 N15918 10
D15918 N15918 0 diode
R15919 N15918 N15919 10
D15919 N15919 0 diode
R15920 N15919 N15920 10
D15920 N15920 0 diode
R15921 N15920 N15921 10
D15921 N15921 0 diode
R15922 N15921 N15922 10
D15922 N15922 0 diode
R15923 N15922 N15923 10
D15923 N15923 0 diode
R15924 N15923 N15924 10
D15924 N15924 0 diode
R15925 N15924 N15925 10
D15925 N15925 0 diode
R15926 N15925 N15926 10
D15926 N15926 0 diode
R15927 N15926 N15927 10
D15927 N15927 0 diode
R15928 N15927 N15928 10
D15928 N15928 0 diode
R15929 N15928 N15929 10
D15929 N15929 0 diode
R15930 N15929 N15930 10
D15930 N15930 0 diode
R15931 N15930 N15931 10
D15931 N15931 0 diode
R15932 N15931 N15932 10
D15932 N15932 0 diode
R15933 N15932 N15933 10
D15933 N15933 0 diode
R15934 N15933 N15934 10
D15934 N15934 0 diode
R15935 N15934 N15935 10
D15935 N15935 0 diode
R15936 N15935 N15936 10
D15936 N15936 0 diode
R15937 N15936 N15937 10
D15937 N15937 0 diode
R15938 N15937 N15938 10
D15938 N15938 0 diode
R15939 N15938 N15939 10
D15939 N15939 0 diode
R15940 N15939 N15940 10
D15940 N15940 0 diode
R15941 N15940 N15941 10
D15941 N15941 0 diode
R15942 N15941 N15942 10
D15942 N15942 0 diode
R15943 N15942 N15943 10
D15943 N15943 0 diode
R15944 N15943 N15944 10
D15944 N15944 0 diode
R15945 N15944 N15945 10
D15945 N15945 0 diode
R15946 N15945 N15946 10
D15946 N15946 0 diode
R15947 N15946 N15947 10
D15947 N15947 0 diode
R15948 N15947 N15948 10
D15948 N15948 0 diode
R15949 N15948 N15949 10
D15949 N15949 0 diode
R15950 N15949 N15950 10
D15950 N15950 0 diode
R15951 N15950 N15951 10
D15951 N15951 0 diode
R15952 N15951 N15952 10
D15952 N15952 0 diode
R15953 N15952 N15953 10
D15953 N15953 0 diode
R15954 N15953 N15954 10
D15954 N15954 0 diode
R15955 N15954 N15955 10
D15955 N15955 0 diode
R15956 N15955 N15956 10
D15956 N15956 0 diode
R15957 N15956 N15957 10
D15957 N15957 0 diode
R15958 N15957 N15958 10
D15958 N15958 0 diode
R15959 N15958 N15959 10
D15959 N15959 0 diode
R15960 N15959 N15960 10
D15960 N15960 0 diode
R15961 N15960 N15961 10
D15961 N15961 0 diode
R15962 N15961 N15962 10
D15962 N15962 0 diode
R15963 N15962 N15963 10
D15963 N15963 0 diode
R15964 N15963 N15964 10
D15964 N15964 0 diode
R15965 N15964 N15965 10
D15965 N15965 0 diode
R15966 N15965 N15966 10
D15966 N15966 0 diode
R15967 N15966 N15967 10
D15967 N15967 0 diode
R15968 N15967 N15968 10
D15968 N15968 0 diode
R15969 N15968 N15969 10
D15969 N15969 0 diode
R15970 N15969 N15970 10
D15970 N15970 0 diode
R15971 N15970 N15971 10
D15971 N15971 0 diode
R15972 N15971 N15972 10
D15972 N15972 0 diode
R15973 N15972 N15973 10
D15973 N15973 0 diode
R15974 N15973 N15974 10
D15974 N15974 0 diode
R15975 N15974 N15975 10
D15975 N15975 0 diode
R15976 N15975 N15976 10
D15976 N15976 0 diode
R15977 N15976 N15977 10
D15977 N15977 0 diode
R15978 N15977 N15978 10
D15978 N15978 0 diode
R15979 N15978 N15979 10
D15979 N15979 0 diode
R15980 N15979 N15980 10
D15980 N15980 0 diode
R15981 N15980 N15981 10
D15981 N15981 0 diode
R15982 N15981 N15982 10
D15982 N15982 0 diode
R15983 N15982 N15983 10
D15983 N15983 0 diode
R15984 N15983 N15984 10
D15984 N15984 0 diode
R15985 N15984 N15985 10
D15985 N15985 0 diode
R15986 N15985 N15986 10
D15986 N15986 0 diode
R15987 N15986 N15987 10
D15987 N15987 0 diode
R15988 N15987 N15988 10
D15988 N15988 0 diode
R15989 N15988 N15989 10
D15989 N15989 0 diode
R15990 N15989 N15990 10
D15990 N15990 0 diode
R15991 N15990 N15991 10
D15991 N15991 0 diode
R15992 N15991 N15992 10
D15992 N15992 0 diode
R15993 N15992 N15993 10
D15993 N15993 0 diode
R15994 N15993 N15994 10
D15994 N15994 0 diode
R15995 N15994 N15995 10
D15995 N15995 0 diode
R15996 N15995 N15996 10
D15996 N15996 0 diode
R15997 N15996 N15997 10
D15997 N15997 0 diode
R15998 N15997 N15998 10
D15998 N15998 0 diode
R15999 N15998 N15999 10
D15999 N15999 0 diode
R16000 N15999 N16000 10
D16000 N16000 0 diode
R16001 N16000 N16001 10
D16001 N16001 0 diode
R16002 N16001 N16002 10
D16002 N16002 0 diode
R16003 N16002 N16003 10
D16003 N16003 0 diode
R16004 N16003 N16004 10
D16004 N16004 0 diode
R16005 N16004 N16005 10
D16005 N16005 0 diode
R16006 N16005 N16006 10
D16006 N16006 0 diode
R16007 N16006 N16007 10
D16007 N16007 0 diode
R16008 N16007 N16008 10
D16008 N16008 0 diode
R16009 N16008 N16009 10
D16009 N16009 0 diode
R16010 N16009 N16010 10
D16010 N16010 0 diode
R16011 N16010 N16011 10
D16011 N16011 0 diode
R16012 N16011 N16012 10
D16012 N16012 0 diode
R16013 N16012 N16013 10
D16013 N16013 0 diode
R16014 N16013 N16014 10
D16014 N16014 0 diode
R16015 N16014 N16015 10
D16015 N16015 0 diode
R16016 N16015 N16016 10
D16016 N16016 0 diode
R16017 N16016 N16017 10
D16017 N16017 0 diode
R16018 N16017 N16018 10
D16018 N16018 0 diode
R16019 N16018 N16019 10
D16019 N16019 0 diode
R16020 N16019 N16020 10
D16020 N16020 0 diode
R16021 N16020 N16021 10
D16021 N16021 0 diode
R16022 N16021 N16022 10
D16022 N16022 0 diode
R16023 N16022 N16023 10
D16023 N16023 0 diode
R16024 N16023 N16024 10
D16024 N16024 0 diode
R16025 N16024 N16025 10
D16025 N16025 0 diode
R16026 N16025 N16026 10
D16026 N16026 0 diode
R16027 N16026 N16027 10
D16027 N16027 0 diode
R16028 N16027 N16028 10
D16028 N16028 0 diode
R16029 N16028 N16029 10
D16029 N16029 0 diode
R16030 N16029 N16030 10
D16030 N16030 0 diode
R16031 N16030 N16031 10
D16031 N16031 0 diode
R16032 N16031 N16032 10
D16032 N16032 0 diode
R16033 N16032 N16033 10
D16033 N16033 0 diode
R16034 N16033 N16034 10
D16034 N16034 0 diode
R16035 N16034 N16035 10
D16035 N16035 0 diode
R16036 N16035 N16036 10
D16036 N16036 0 diode
R16037 N16036 N16037 10
D16037 N16037 0 diode
R16038 N16037 N16038 10
D16038 N16038 0 diode
R16039 N16038 N16039 10
D16039 N16039 0 diode
R16040 N16039 N16040 10
D16040 N16040 0 diode
R16041 N16040 N16041 10
D16041 N16041 0 diode
R16042 N16041 N16042 10
D16042 N16042 0 diode
R16043 N16042 N16043 10
D16043 N16043 0 diode
R16044 N16043 N16044 10
D16044 N16044 0 diode
R16045 N16044 N16045 10
D16045 N16045 0 diode
R16046 N16045 N16046 10
D16046 N16046 0 diode
R16047 N16046 N16047 10
D16047 N16047 0 diode
R16048 N16047 N16048 10
D16048 N16048 0 diode
R16049 N16048 N16049 10
D16049 N16049 0 diode
R16050 N16049 N16050 10
D16050 N16050 0 diode
R16051 N16050 N16051 10
D16051 N16051 0 diode
R16052 N16051 N16052 10
D16052 N16052 0 diode
R16053 N16052 N16053 10
D16053 N16053 0 diode
R16054 N16053 N16054 10
D16054 N16054 0 diode
R16055 N16054 N16055 10
D16055 N16055 0 diode
R16056 N16055 N16056 10
D16056 N16056 0 diode
R16057 N16056 N16057 10
D16057 N16057 0 diode
R16058 N16057 N16058 10
D16058 N16058 0 diode
R16059 N16058 N16059 10
D16059 N16059 0 diode
R16060 N16059 N16060 10
D16060 N16060 0 diode
R16061 N16060 N16061 10
D16061 N16061 0 diode
R16062 N16061 N16062 10
D16062 N16062 0 diode
R16063 N16062 N16063 10
D16063 N16063 0 diode
R16064 N16063 N16064 10
D16064 N16064 0 diode
R16065 N16064 N16065 10
D16065 N16065 0 diode
R16066 N16065 N16066 10
D16066 N16066 0 diode
R16067 N16066 N16067 10
D16067 N16067 0 diode
R16068 N16067 N16068 10
D16068 N16068 0 diode
R16069 N16068 N16069 10
D16069 N16069 0 diode
R16070 N16069 N16070 10
D16070 N16070 0 diode
R16071 N16070 N16071 10
D16071 N16071 0 diode
R16072 N16071 N16072 10
D16072 N16072 0 diode
R16073 N16072 N16073 10
D16073 N16073 0 diode
R16074 N16073 N16074 10
D16074 N16074 0 diode
R16075 N16074 N16075 10
D16075 N16075 0 diode
R16076 N16075 N16076 10
D16076 N16076 0 diode
R16077 N16076 N16077 10
D16077 N16077 0 diode
R16078 N16077 N16078 10
D16078 N16078 0 diode
R16079 N16078 N16079 10
D16079 N16079 0 diode
R16080 N16079 N16080 10
D16080 N16080 0 diode
R16081 N16080 N16081 10
D16081 N16081 0 diode
R16082 N16081 N16082 10
D16082 N16082 0 diode
R16083 N16082 N16083 10
D16083 N16083 0 diode
R16084 N16083 N16084 10
D16084 N16084 0 diode
R16085 N16084 N16085 10
D16085 N16085 0 diode
R16086 N16085 N16086 10
D16086 N16086 0 diode
R16087 N16086 N16087 10
D16087 N16087 0 diode
R16088 N16087 N16088 10
D16088 N16088 0 diode
R16089 N16088 N16089 10
D16089 N16089 0 diode
R16090 N16089 N16090 10
D16090 N16090 0 diode
R16091 N16090 N16091 10
D16091 N16091 0 diode
R16092 N16091 N16092 10
D16092 N16092 0 diode
R16093 N16092 N16093 10
D16093 N16093 0 diode
R16094 N16093 N16094 10
D16094 N16094 0 diode
R16095 N16094 N16095 10
D16095 N16095 0 diode
R16096 N16095 N16096 10
D16096 N16096 0 diode
R16097 N16096 N16097 10
D16097 N16097 0 diode
R16098 N16097 N16098 10
D16098 N16098 0 diode
R16099 N16098 N16099 10
D16099 N16099 0 diode
R16100 N16099 N16100 10
D16100 N16100 0 diode
R16101 N16100 N16101 10
D16101 N16101 0 diode
R16102 N16101 N16102 10
D16102 N16102 0 diode
R16103 N16102 N16103 10
D16103 N16103 0 diode
R16104 N16103 N16104 10
D16104 N16104 0 diode
R16105 N16104 N16105 10
D16105 N16105 0 diode
R16106 N16105 N16106 10
D16106 N16106 0 diode
R16107 N16106 N16107 10
D16107 N16107 0 diode
R16108 N16107 N16108 10
D16108 N16108 0 diode
R16109 N16108 N16109 10
D16109 N16109 0 diode
R16110 N16109 N16110 10
D16110 N16110 0 diode
R16111 N16110 N16111 10
D16111 N16111 0 diode
R16112 N16111 N16112 10
D16112 N16112 0 diode
R16113 N16112 N16113 10
D16113 N16113 0 diode
R16114 N16113 N16114 10
D16114 N16114 0 diode
R16115 N16114 N16115 10
D16115 N16115 0 diode
R16116 N16115 N16116 10
D16116 N16116 0 diode
R16117 N16116 N16117 10
D16117 N16117 0 diode
R16118 N16117 N16118 10
D16118 N16118 0 diode
R16119 N16118 N16119 10
D16119 N16119 0 diode
R16120 N16119 N16120 10
D16120 N16120 0 diode
R16121 N16120 N16121 10
D16121 N16121 0 diode
R16122 N16121 N16122 10
D16122 N16122 0 diode
R16123 N16122 N16123 10
D16123 N16123 0 diode
R16124 N16123 N16124 10
D16124 N16124 0 diode
R16125 N16124 N16125 10
D16125 N16125 0 diode
R16126 N16125 N16126 10
D16126 N16126 0 diode
R16127 N16126 N16127 10
D16127 N16127 0 diode
R16128 N16127 N16128 10
D16128 N16128 0 diode
R16129 N16128 N16129 10
D16129 N16129 0 diode
R16130 N16129 N16130 10
D16130 N16130 0 diode
R16131 N16130 N16131 10
D16131 N16131 0 diode
R16132 N16131 N16132 10
D16132 N16132 0 diode
R16133 N16132 N16133 10
D16133 N16133 0 diode
R16134 N16133 N16134 10
D16134 N16134 0 diode
R16135 N16134 N16135 10
D16135 N16135 0 diode
R16136 N16135 N16136 10
D16136 N16136 0 diode
R16137 N16136 N16137 10
D16137 N16137 0 diode
R16138 N16137 N16138 10
D16138 N16138 0 diode
R16139 N16138 N16139 10
D16139 N16139 0 diode
R16140 N16139 N16140 10
D16140 N16140 0 diode
R16141 N16140 N16141 10
D16141 N16141 0 diode
R16142 N16141 N16142 10
D16142 N16142 0 diode
R16143 N16142 N16143 10
D16143 N16143 0 diode
R16144 N16143 N16144 10
D16144 N16144 0 diode
R16145 N16144 N16145 10
D16145 N16145 0 diode
R16146 N16145 N16146 10
D16146 N16146 0 diode
R16147 N16146 N16147 10
D16147 N16147 0 diode
R16148 N16147 N16148 10
D16148 N16148 0 diode
R16149 N16148 N16149 10
D16149 N16149 0 diode
R16150 N16149 N16150 10
D16150 N16150 0 diode
R16151 N16150 N16151 10
D16151 N16151 0 diode
R16152 N16151 N16152 10
D16152 N16152 0 diode
R16153 N16152 N16153 10
D16153 N16153 0 diode
R16154 N16153 N16154 10
D16154 N16154 0 diode
R16155 N16154 N16155 10
D16155 N16155 0 diode
R16156 N16155 N16156 10
D16156 N16156 0 diode
R16157 N16156 N16157 10
D16157 N16157 0 diode
R16158 N16157 N16158 10
D16158 N16158 0 diode
R16159 N16158 N16159 10
D16159 N16159 0 diode
R16160 N16159 N16160 10
D16160 N16160 0 diode
R16161 N16160 N16161 10
D16161 N16161 0 diode
R16162 N16161 N16162 10
D16162 N16162 0 diode
R16163 N16162 N16163 10
D16163 N16163 0 diode
R16164 N16163 N16164 10
D16164 N16164 0 diode
R16165 N16164 N16165 10
D16165 N16165 0 diode
R16166 N16165 N16166 10
D16166 N16166 0 diode
R16167 N16166 N16167 10
D16167 N16167 0 diode
R16168 N16167 N16168 10
D16168 N16168 0 diode
R16169 N16168 N16169 10
D16169 N16169 0 diode
R16170 N16169 N16170 10
D16170 N16170 0 diode
R16171 N16170 N16171 10
D16171 N16171 0 diode
R16172 N16171 N16172 10
D16172 N16172 0 diode
R16173 N16172 N16173 10
D16173 N16173 0 diode
R16174 N16173 N16174 10
D16174 N16174 0 diode
R16175 N16174 N16175 10
D16175 N16175 0 diode
R16176 N16175 N16176 10
D16176 N16176 0 diode
R16177 N16176 N16177 10
D16177 N16177 0 diode
R16178 N16177 N16178 10
D16178 N16178 0 diode
R16179 N16178 N16179 10
D16179 N16179 0 diode
R16180 N16179 N16180 10
D16180 N16180 0 diode
R16181 N16180 N16181 10
D16181 N16181 0 diode
R16182 N16181 N16182 10
D16182 N16182 0 diode
R16183 N16182 N16183 10
D16183 N16183 0 diode
R16184 N16183 N16184 10
D16184 N16184 0 diode
R16185 N16184 N16185 10
D16185 N16185 0 diode
R16186 N16185 N16186 10
D16186 N16186 0 diode
R16187 N16186 N16187 10
D16187 N16187 0 diode
R16188 N16187 N16188 10
D16188 N16188 0 diode
R16189 N16188 N16189 10
D16189 N16189 0 diode
R16190 N16189 N16190 10
D16190 N16190 0 diode
R16191 N16190 N16191 10
D16191 N16191 0 diode
R16192 N16191 N16192 10
D16192 N16192 0 diode
R16193 N16192 N16193 10
D16193 N16193 0 diode
R16194 N16193 N16194 10
D16194 N16194 0 diode
R16195 N16194 N16195 10
D16195 N16195 0 diode
R16196 N16195 N16196 10
D16196 N16196 0 diode
R16197 N16196 N16197 10
D16197 N16197 0 diode
R16198 N16197 N16198 10
D16198 N16198 0 diode
R16199 N16198 N16199 10
D16199 N16199 0 diode
R16200 N16199 N16200 10
D16200 N16200 0 diode
R16201 N16200 N16201 10
D16201 N16201 0 diode
R16202 N16201 N16202 10
D16202 N16202 0 diode
R16203 N16202 N16203 10
D16203 N16203 0 diode
R16204 N16203 N16204 10
D16204 N16204 0 diode
R16205 N16204 N16205 10
D16205 N16205 0 diode
R16206 N16205 N16206 10
D16206 N16206 0 diode
R16207 N16206 N16207 10
D16207 N16207 0 diode
R16208 N16207 N16208 10
D16208 N16208 0 diode
R16209 N16208 N16209 10
D16209 N16209 0 diode
R16210 N16209 N16210 10
D16210 N16210 0 diode
R16211 N16210 N16211 10
D16211 N16211 0 diode
R16212 N16211 N16212 10
D16212 N16212 0 diode
R16213 N16212 N16213 10
D16213 N16213 0 diode
R16214 N16213 N16214 10
D16214 N16214 0 diode
R16215 N16214 N16215 10
D16215 N16215 0 diode
R16216 N16215 N16216 10
D16216 N16216 0 diode
R16217 N16216 N16217 10
D16217 N16217 0 diode
R16218 N16217 N16218 10
D16218 N16218 0 diode
R16219 N16218 N16219 10
D16219 N16219 0 diode
R16220 N16219 N16220 10
D16220 N16220 0 diode
R16221 N16220 N16221 10
D16221 N16221 0 diode
R16222 N16221 N16222 10
D16222 N16222 0 diode
R16223 N16222 N16223 10
D16223 N16223 0 diode
R16224 N16223 N16224 10
D16224 N16224 0 diode
R16225 N16224 N16225 10
D16225 N16225 0 diode
R16226 N16225 N16226 10
D16226 N16226 0 diode
R16227 N16226 N16227 10
D16227 N16227 0 diode
R16228 N16227 N16228 10
D16228 N16228 0 diode
R16229 N16228 N16229 10
D16229 N16229 0 diode
R16230 N16229 N16230 10
D16230 N16230 0 diode
R16231 N16230 N16231 10
D16231 N16231 0 diode
R16232 N16231 N16232 10
D16232 N16232 0 diode
R16233 N16232 N16233 10
D16233 N16233 0 diode
R16234 N16233 N16234 10
D16234 N16234 0 diode
R16235 N16234 N16235 10
D16235 N16235 0 diode
R16236 N16235 N16236 10
D16236 N16236 0 diode
R16237 N16236 N16237 10
D16237 N16237 0 diode
R16238 N16237 N16238 10
D16238 N16238 0 diode
R16239 N16238 N16239 10
D16239 N16239 0 diode
R16240 N16239 N16240 10
D16240 N16240 0 diode
R16241 N16240 N16241 10
D16241 N16241 0 diode
R16242 N16241 N16242 10
D16242 N16242 0 diode
R16243 N16242 N16243 10
D16243 N16243 0 diode
R16244 N16243 N16244 10
D16244 N16244 0 diode
R16245 N16244 N16245 10
D16245 N16245 0 diode
R16246 N16245 N16246 10
D16246 N16246 0 diode
R16247 N16246 N16247 10
D16247 N16247 0 diode
R16248 N16247 N16248 10
D16248 N16248 0 diode
R16249 N16248 N16249 10
D16249 N16249 0 diode
R16250 N16249 N16250 10
D16250 N16250 0 diode
R16251 N16250 N16251 10
D16251 N16251 0 diode
R16252 N16251 N16252 10
D16252 N16252 0 diode
R16253 N16252 N16253 10
D16253 N16253 0 diode
R16254 N16253 N16254 10
D16254 N16254 0 diode
R16255 N16254 N16255 10
D16255 N16255 0 diode
R16256 N16255 N16256 10
D16256 N16256 0 diode
R16257 N16256 N16257 10
D16257 N16257 0 diode
R16258 N16257 N16258 10
D16258 N16258 0 diode
R16259 N16258 N16259 10
D16259 N16259 0 diode
R16260 N16259 N16260 10
D16260 N16260 0 diode
R16261 N16260 N16261 10
D16261 N16261 0 diode
R16262 N16261 N16262 10
D16262 N16262 0 diode
R16263 N16262 N16263 10
D16263 N16263 0 diode
R16264 N16263 N16264 10
D16264 N16264 0 diode
R16265 N16264 N16265 10
D16265 N16265 0 diode
R16266 N16265 N16266 10
D16266 N16266 0 diode
R16267 N16266 N16267 10
D16267 N16267 0 diode
R16268 N16267 N16268 10
D16268 N16268 0 diode
R16269 N16268 N16269 10
D16269 N16269 0 diode
R16270 N16269 N16270 10
D16270 N16270 0 diode
R16271 N16270 N16271 10
D16271 N16271 0 diode
R16272 N16271 N16272 10
D16272 N16272 0 diode
R16273 N16272 N16273 10
D16273 N16273 0 diode
R16274 N16273 N16274 10
D16274 N16274 0 diode
R16275 N16274 N16275 10
D16275 N16275 0 diode
R16276 N16275 N16276 10
D16276 N16276 0 diode
R16277 N16276 N16277 10
D16277 N16277 0 diode
R16278 N16277 N16278 10
D16278 N16278 0 diode
R16279 N16278 N16279 10
D16279 N16279 0 diode
R16280 N16279 N16280 10
D16280 N16280 0 diode
R16281 N16280 N16281 10
D16281 N16281 0 diode
R16282 N16281 N16282 10
D16282 N16282 0 diode
R16283 N16282 N16283 10
D16283 N16283 0 diode
R16284 N16283 N16284 10
D16284 N16284 0 diode
R16285 N16284 N16285 10
D16285 N16285 0 diode
R16286 N16285 N16286 10
D16286 N16286 0 diode
R16287 N16286 N16287 10
D16287 N16287 0 diode
R16288 N16287 N16288 10
D16288 N16288 0 diode
R16289 N16288 N16289 10
D16289 N16289 0 diode
R16290 N16289 N16290 10
D16290 N16290 0 diode
R16291 N16290 N16291 10
D16291 N16291 0 diode
R16292 N16291 N16292 10
D16292 N16292 0 diode
R16293 N16292 N16293 10
D16293 N16293 0 diode
R16294 N16293 N16294 10
D16294 N16294 0 diode
R16295 N16294 N16295 10
D16295 N16295 0 diode
R16296 N16295 N16296 10
D16296 N16296 0 diode
R16297 N16296 N16297 10
D16297 N16297 0 diode
R16298 N16297 N16298 10
D16298 N16298 0 diode
R16299 N16298 N16299 10
D16299 N16299 0 diode
R16300 N16299 N16300 10
D16300 N16300 0 diode
R16301 N16300 N16301 10
D16301 N16301 0 diode
R16302 N16301 N16302 10
D16302 N16302 0 diode
R16303 N16302 N16303 10
D16303 N16303 0 diode
R16304 N16303 N16304 10
D16304 N16304 0 diode
R16305 N16304 N16305 10
D16305 N16305 0 diode
R16306 N16305 N16306 10
D16306 N16306 0 diode
R16307 N16306 N16307 10
D16307 N16307 0 diode
R16308 N16307 N16308 10
D16308 N16308 0 diode
R16309 N16308 N16309 10
D16309 N16309 0 diode
R16310 N16309 N16310 10
D16310 N16310 0 diode
R16311 N16310 N16311 10
D16311 N16311 0 diode
R16312 N16311 N16312 10
D16312 N16312 0 diode
R16313 N16312 N16313 10
D16313 N16313 0 diode
R16314 N16313 N16314 10
D16314 N16314 0 diode
R16315 N16314 N16315 10
D16315 N16315 0 diode
R16316 N16315 N16316 10
D16316 N16316 0 diode
R16317 N16316 N16317 10
D16317 N16317 0 diode
R16318 N16317 N16318 10
D16318 N16318 0 diode
R16319 N16318 N16319 10
D16319 N16319 0 diode
R16320 N16319 N16320 10
D16320 N16320 0 diode
R16321 N16320 N16321 10
D16321 N16321 0 diode
R16322 N16321 N16322 10
D16322 N16322 0 diode
R16323 N16322 N16323 10
D16323 N16323 0 diode
R16324 N16323 N16324 10
D16324 N16324 0 diode
R16325 N16324 N16325 10
D16325 N16325 0 diode
R16326 N16325 N16326 10
D16326 N16326 0 diode
R16327 N16326 N16327 10
D16327 N16327 0 diode
R16328 N16327 N16328 10
D16328 N16328 0 diode
R16329 N16328 N16329 10
D16329 N16329 0 diode
R16330 N16329 N16330 10
D16330 N16330 0 diode
R16331 N16330 N16331 10
D16331 N16331 0 diode
R16332 N16331 N16332 10
D16332 N16332 0 diode
R16333 N16332 N16333 10
D16333 N16333 0 diode
R16334 N16333 N16334 10
D16334 N16334 0 diode
R16335 N16334 N16335 10
D16335 N16335 0 diode
R16336 N16335 N16336 10
D16336 N16336 0 diode
R16337 N16336 N16337 10
D16337 N16337 0 diode
R16338 N16337 N16338 10
D16338 N16338 0 diode
R16339 N16338 N16339 10
D16339 N16339 0 diode
R16340 N16339 N16340 10
D16340 N16340 0 diode
R16341 N16340 N16341 10
D16341 N16341 0 diode
R16342 N16341 N16342 10
D16342 N16342 0 diode
R16343 N16342 N16343 10
D16343 N16343 0 diode
R16344 N16343 N16344 10
D16344 N16344 0 diode
R16345 N16344 N16345 10
D16345 N16345 0 diode
R16346 N16345 N16346 10
D16346 N16346 0 diode
R16347 N16346 N16347 10
D16347 N16347 0 diode
R16348 N16347 N16348 10
D16348 N16348 0 diode
R16349 N16348 N16349 10
D16349 N16349 0 diode
R16350 N16349 N16350 10
D16350 N16350 0 diode
R16351 N16350 N16351 10
D16351 N16351 0 diode
R16352 N16351 N16352 10
D16352 N16352 0 diode
R16353 N16352 N16353 10
D16353 N16353 0 diode
R16354 N16353 N16354 10
D16354 N16354 0 diode
R16355 N16354 N16355 10
D16355 N16355 0 diode
R16356 N16355 N16356 10
D16356 N16356 0 diode
R16357 N16356 N16357 10
D16357 N16357 0 diode
R16358 N16357 N16358 10
D16358 N16358 0 diode
R16359 N16358 N16359 10
D16359 N16359 0 diode
R16360 N16359 N16360 10
D16360 N16360 0 diode
R16361 N16360 N16361 10
D16361 N16361 0 diode
R16362 N16361 N16362 10
D16362 N16362 0 diode
R16363 N16362 N16363 10
D16363 N16363 0 diode
R16364 N16363 N16364 10
D16364 N16364 0 diode
R16365 N16364 N16365 10
D16365 N16365 0 diode
R16366 N16365 N16366 10
D16366 N16366 0 diode
R16367 N16366 N16367 10
D16367 N16367 0 diode
R16368 N16367 N16368 10
D16368 N16368 0 diode
R16369 N16368 N16369 10
D16369 N16369 0 diode
R16370 N16369 N16370 10
D16370 N16370 0 diode
R16371 N16370 N16371 10
D16371 N16371 0 diode
R16372 N16371 N16372 10
D16372 N16372 0 diode
R16373 N16372 N16373 10
D16373 N16373 0 diode
R16374 N16373 N16374 10
D16374 N16374 0 diode
R16375 N16374 N16375 10
D16375 N16375 0 diode
R16376 N16375 N16376 10
D16376 N16376 0 diode
R16377 N16376 N16377 10
D16377 N16377 0 diode
R16378 N16377 N16378 10
D16378 N16378 0 diode
R16379 N16378 N16379 10
D16379 N16379 0 diode
R16380 N16379 N16380 10
D16380 N16380 0 diode
R16381 N16380 N16381 10
D16381 N16381 0 diode
R16382 N16381 N16382 10
D16382 N16382 0 diode
R16383 N16382 N16383 10
D16383 N16383 0 diode
R16384 N16383 N16384 10
D16384 N16384 0 diode
R16385 N16384 N16385 10
D16385 N16385 0 diode
R16386 N16385 N16386 10
D16386 N16386 0 diode
R16387 N16386 N16387 10
D16387 N16387 0 diode
R16388 N16387 N16388 10
D16388 N16388 0 diode
R16389 N16388 N16389 10
D16389 N16389 0 diode
R16390 N16389 N16390 10
D16390 N16390 0 diode
R16391 N16390 N16391 10
D16391 N16391 0 diode
R16392 N16391 N16392 10
D16392 N16392 0 diode
R16393 N16392 N16393 10
D16393 N16393 0 diode
R16394 N16393 N16394 10
D16394 N16394 0 diode
R16395 N16394 N16395 10
D16395 N16395 0 diode
R16396 N16395 N16396 10
D16396 N16396 0 diode
R16397 N16396 N16397 10
D16397 N16397 0 diode
R16398 N16397 N16398 10
D16398 N16398 0 diode
R16399 N16398 N16399 10
D16399 N16399 0 diode
R16400 N16399 N16400 10
D16400 N16400 0 diode
R16401 N16400 N16401 10
D16401 N16401 0 diode
R16402 N16401 N16402 10
D16402 N16402 0 diode
R16403 N16402 N16403 10
D16403 N16403 0 diode
R16404 N16403 N16404 10
D16404 N16404 0 diode
R16405 N16404 N16405 10
D16405 N16405 0 diode
R16406 N16405 N16406 10
D16406 N16406 0 diode
R16407 N16406 N16407 10
D16407 N16407 0 diode
R16408 N16407 N16408 10
D16408 N16408 0 diode
R16409 N16408 N16409 10
D16409 N16409 0 diode
R16410 N16409 N16410 10
D16410 N16410 0 diode
R16411 N16410 N16411 10
D16411 N16411 0 diode
R16412 N16411 N16412 10
D16412 N16412 0 diode
R16413 N16412 N16413 10
D16413 N16413 0 diode
R16414 N16413 N16414 10
D16414 N16414 0 diode
R16415 N16414 N16415 10
D16415 N16415 0 diode
R16416 N16415 N16416 10
D16416 N16416 0 diode
R16417 N16416 N16417 10
D16417 N16417 0 diode
R16418 N16417 N16418 10
D16418 N16418 0 diode
R16419 N16418 N16419 10
D16419 N16419 0 diode
R16420 N16419 N16420 10
D16420 N16420 0 diode
R16421 N16420 N16421 10
D16421 N16421 0 diode
R16422 N16421 N16422 10
D16422 N16422 0 diode
R16423 N16422 N16423 10
D16423 N16423 0 diode
R16424 N16423 N16424 10
D16424 N16424 0 diode
R16425 N16424 N16425 10
D16425 N16425 0 diode
R16426 N16425 N16426 10
D16426 N16426 0 diode
R16427 N16426 N16427 10
D16427 N16427 0 diode
R16428 N16427 N16428 10
D16428 N16428 0 diode
R16429 N16428 N16429 10
D16429 N16429 0 diode
R16430 N16429 N16430 10
D16430 N16430 0 diode
R16431 N16430 N16431 10
D16431 N16431 0 diode
R16432 N16431 N16432 10
D16432 N16432 0 diode
R16433 N16432 N16433 10
D16433 N16433 0 diode
R16434 N16433 N16434 10
D16434 N16434 0 diode
R16435 N16434 N16435 10
D16435 N16435 0 diode
R16436 N16435 N16436 10
D16436 N16436 0 diode
R16437 N16436 N16437 10
D16437 N16437 0 diode
R16438 N16437 N16438 10
D16438 N16438 0 diode
R16439 N16438 N16439 10
D16439 N16439 0 diode
R16440 N16439 N16440 10
D16440 N16440 0 diode
R16441 N16440 N16441 10
D16441 N16441 0 diode
R16442 N16441 N16442 10
D16442 N16442 0 diode
R16443 N16442 N16443 10
D16443 N16443 0 diode
R16444 N16443 N16444 10
D16444 N16444 0 diode
R16445 N16444 N16445 10
D16445 N16445 0 diode
R16446 N16445 N16446 10
D16446 N16446 0 diode
R16447 N16446 N16447 10
D16447 N16447 0 diode
R16448 N16447 N16448 10
D16448 N16448 0 diode
R16449 N16448 N16449 10
D16449 N16449 0 diode
R16450 N16449 N16450 10
D16450 N16450 0 diode
R16451 N16450 N16451 10
D16451 N16451 0 diode
R16452 N16451 N16452 10
D16452 N16452 0 diode
R16453 N16452 N16453 10
D16453 N16453 0 diode
R16454 N16453 N16454 10
D16454 N16454 0 diode
R16455 N16454 N16455 10
D16455 N16455 0 diode
R16456 N16455 N16456 10
D16456 N16456 0 diode
R16457 N16456 N16457 10
D16457 N16457 0 diode
R16458 N16457 N16458 10
D16458 N16458 0 diode
R16459 N16458 N16459 10
D16459 N16459 0 diode
R16460 N16459 N16460 10
D16460 N16460 0 diode
R16461 N16460 N16461 10
D16461 N16461 0 diode
R16462 N16461 N16462 10
D16462 N16462 0 diode
R16463 N16462 N16463 10
D16463 N16463 0 diode
R16464 N16463 N16464 10
D16464 N16464 0 diode
R16465 N16464 N16465 10
D16465 N16465 0 diode
R16466 N16465 N16466 10
D16466 N16466 0 diode
R16467 N16466 N16467 10
D16467 N16467 0 diode
R16468 N16467 N16468 10
D16468 N16468 0 diode
R16469 N16468 N16469 10
D16469 N16469 0 diode
R16470 N16469 N16470 10
D16470 N16470 0 diode
R16471 N16470 N16471 10
D16471 N16471 0 diode
R16472 N16471 N16472 10
D16472 N16472 0 diode
R16473 N16472 N16473 10
D16473 N16473 0 diode
R16474 N16473 N16474 10
D16474 N16474 0 diode
R16475 N16474 N16475 10
D16475 N16475 0 diode
R16476 N16475 N16476 10
D16476 N16476 0 diode
R16477 N16476 N16477 10
D16477 N16477 0 diode
R16478 N16477 N16478 10
D16478 N16478 0 diode
R16479 N16478 N16479 10
D16479 N16479 0 diode
R16480 N16479 N16480 10
D16480 N16480 0 diode
R16481 N16480 N16481 10
D16481 N16481 0 diode
R16482 N16481 N16482 10
D16482 N16482 0 diode
R16483 N16482 N16483 10
D16483 N16483 0 diode
R16484 N16483 N16484 10
D16484 N16484 0 diode
R16485 N16484 N16485 10
D16485 N16485 0 diode
R16486 N16485 N16486 10
D16486 N16486 0 diode
R16487 N16486 N16487 10
D16487 N16487 0 diode
R16488 N16487 N16488 10
D16488 N16488 0 diode
R16489 N16488 N16489 10
D16489 N16489 0 diode
R16490 N16489 N16490 10
D16490 N16490 0 diode
R16491 N16490 N16491 10
D16491 N16491 0 diode
R16492 N16491 N16492 10
D16492 N16492 0 diode
R16493 N16492 N16493 10
D16493 N16493 0 diode
R16494 N16493 N16494 10
D16494 N16494 0 diode
R16495 N16494 N16495 10
D16495 N16495 0 diode
R16496 N16495 N16496 10
D16496 N16496 0 diode
R16497 N16496 N16497 10
D16497 N16497 0 diode
R16498 N16497 N16498 10
D16498 N16498 0 diode
R16499 N16498 N16499 10
D16499 N16499 0 diode
R16500 N16499 N16500 10
D16500 N16500 0 diode
R16501 N16500 N16501 10
D16501 N16501 0 diode
R16502 N16501 N16502 10
D16502 N16502 0 diode
R16503 N16502 N16503 10
D16503 N16503 0 diode
R16504 N16503 N16504 10
D16504 N16504 0 diode
R16505 N16504 N16505 10
D16505 N16505 0 diode
R16506 N16505 N16506 10
D16506 N16506 0 diode
R16507 N16506 N16507 10
D16507 N16507 0 diode
R16508 N16507 N16508 10
D16508 N16508 0 diode
R16509 N16508 N16509 10
D16509 N16509 0 diode
R16510 N16509 N16510 10
D16510 N16510 0 diode
R16511 N16510 N16511 10
D16511 N16511 0 diode
R16512 N16511 N16512 10
D16512 N16512 0 diode
R16513 N16512 N16513 10
D16513 N16513 0 diode
R16514 N16513 N16514 10
D16514 N16514 0 diode
R16515 N16514 N16515 10
D16515 N16515 0 diode
R16516 N16515 N16516 10
D16516 N16516 0 diode
R16517 N16516 N16517 10
D16517 N16517 0 diode
R16518 N16517 N16518 10
D16518 N16518 0 diode
R16519 N16518 N16519 10
D16519 N16519 0 diode
R16520 N16519 N16520 10
D16520 N16520 0 diode
R16521 N16520 N16521 10
D16521 N16521 0 diode
R16522 N16521 N16522 10
D16522 N16522 0 diode
R16523 N16522 N16523 10
D16523 N16523 0 diode
R16524 N16523 N16524 10
D16524 N16524 0 diode
R16525 N16524 N16525 10
D16525 N16525 0 diode
R16526 N16525 N16526 10
D16526 N16526 0 diode
R16527 N16526 N16527 10
D16527 N16527 0 diode
R16528 N16527 N16528 10
D16528 N16528 0 diode
R16529 N16528 N16529 10
D16529 N16529 0 diode
R16530 N16529 N16530 10
D16530 N16530 0 diode
R16531 N16530 N16531 10
D16531 N16531 0 diode
R16532 N16531 N16532 10
D16532 N16532 0 diode
R16533 N16532 N16533 10
D16533 N16533 0 diode
R16534 N16533 N16534 10
D16534 N16534 0 diode
R16535 N16534 N16535 10
D16535 N16535 0 diode
R16536 N16535 N16536 10
D16536 N16536 0 diode
R16537 N16536 N16537 10
D16537 N16537 0 diode
R16538 N16537 N16538 10
D16538 N16538 0 diode
R16539 N16538 N16539 10
D16539 N16539 0 diode
R16540 N16539 N16540 10
D16540 N16540 0 diode
R16541 N16540 N16541 10
D16541 N16541 0 diode
R16542 N16541 N16542 10
D16542 N16542 0 diode
R16543 N16542 N16543 10
D16543 N16543 0 diode
R16544 N16543 N16544 10
D16544 N16544 0 diode
R16545 N16544 N16545 10
D16545 N16545 0 diode
R16546 N16545 N16546 10
D16546 N16546 0 diode
R16547 N16546 N16547 10
D16547 N16547 0 diode
R16548 N16547 N16548 10
D16548 N16548 0 diode
R16549 N16548 N16549 10
D16549 N16549 0 diode
R16550 N16549 N16550 10
D16550 N16550 0 diode
R16551 N16550 N16551 10
D16551 N16551 0 diode
R16552 N16551 N16552 10
D16552 N16552 0 diode
R16553 N16552 N16553 10
D16553 N16553 0 diode
R16554 N16553 N16554 10
D16554 N16554 0 diode
R16555 N16554 N16555 10
D16555 N16555 0 diode
R16556 N16555 N16556 10
D16556 N16556 0 diode
R16557 N16556 N16557 10
D16557 N16557 0 diode
R16558 N16557 N16558 10
D16558 N16558 0 diode
R16559 N16558 N16559 10
D16559 N16559 0 diode
R16560 N16559 N16560 10
D16560 N16560 0 diode
R16561 N16560 N16561 10
D16561 N16561 0 diode
R16562 N16561 N16562 10
D16562 N16562 0 diode
R16563 N16562 N16563 10
D16563 N16563 0 diode
R16564 N16563 N16564 10
D16564 N16564 0 diode
R16565 N16564 N16565 10
D16565 N16565 0 diode
R16566 N16565 N16566 10
D16566 N16566 0 diode
R16567 N16566 N16567 10
D16567 N16567 0 diode
R16568 N16567 N16568 10
D16568 N16568 0 diode
R16569 N16568 N16569 10
D16569 N16569 0 diode
R16570 N16569 N16570 10
D16570 N16570 0 diode
R16571 N16570 N16571 10
D16571 N16571 0 diode
R16572 N16571 N16572 10
D16572 N16572 0 diode
R16573 N16572 N16573 10
D16573 N16573 0 diode
R16574 N16573 N16574 10
D16574 N16574 0 diode
R16575 N16574 N16575 10
D16575 N16575 0 diode
R16576 N16575 N16576 10
D16576 N16576 0 diode
R16577 N16576 N16577 10
D16577 N16577 0 diode
R16578 N16577 N16578 10
D16578 N16578 0 diode
R16579 N16578 N16579 10
D16579 N16579 0 diode
R16580 N16579 N16580 10
D16580 N16580 0 diode
R16581 N16580 N16581 10
D16581 N16581 0 diode
R16582 N16581 N16582 10
D16582 N16582 0 diode
R16583 N16582 N16583 10
D16583 N16583 0 diode
R16584 N16583 N16584 10
D16584 N16584 0 diode
R16585 N16584 N16585 10
D16585 N16585 0 diode
R16586 N16585 N16586 10
D16586 N16586 0 diode
R16587 N16586 N16587 10
D16587 N16587 0 diode
R16588 N16587 N16588 10
D16588 N16588 0 diode
R16589 N16588 N16589 10
D16589 N16589 0 diode
R16590 N16589 N16590 10
D16590 N16590 0 diode
R16591 N16590 N16591 10
D16591 N16591 0 diode
R16592 N16591 N16592 10
D16592 N16592 0 diode
R16593 N16592 N16593 10
D16593 N16593 0 diode
R16594 N16593 N16594 10
D16594 N16594 0 diode
R16595 N16594 N16595 10
D16595 N16595 0 diode
R16596 N16595 N16596 10
D16596 N16596 0 diode
R16597 N16596 N16597 10
D16597 N16597 0 diode
R16598 N16597 N16598 10
D16598 N16598 0 diode
R16599 N16598 N16599 10
D16599 N16599 0 diode
R16600 N16599 N16600 10
D16600 N16600 0 diode
R16601 N16600 N16601 10
D16601 N16601 0 diode
R16602 N16601 N16602 10
D16602 N16602 0 diode
R16603 N16602 N16603 10
D16603 N16603 0 diode
R16604 N16603 N16604 10
D16604 N16604 0 diode
R16605 N16604 N16605 10
D16605 N16605 0 diode
R16606 N16605 N16606 10
D16606 N16606 0 diode
R16607 N16606 N16607 10
D16607 N16607 0 diode
R16608 N16607 N16608 10
D16608 N16608 0 diode
R16609 N16608 N16609 10
D16609 N16609 0 diode
R16610 N16609 N16610 10
D16610 N16610 0 diode
R16611 N16610 N16611 10
D16611 N16611 0 diode
R16612 N16611 N16612 10
D16612 N16612 0 diode
R16613 N16612 N16613 10
D16613 N16613 0 diode
R16614 N16613 N16614 10
D16614 N16614 0 diode
R16615 N16614 N16615 10
D16615 N16615 0 diode
R16616 N16615 N16616 10
D16616 N16616 0 diode
R16617 N16616 N16617 10
D16617 N16617 0 diode
R16618 N16617 N16618 10
D16618 N16618 0 diode
R16619 N16618 N16619 10
D16619 N16619 0 diode
R16620 N16619 N16620 10
D16620 N16620 0 diode
R16621 N16620 N16621 10
D16621 N16621 0 diode
R16622 N16621 N16622 10
D16622 N16622 0 diode
R16623 N16622 N16623 10
D16623 N16623 0 diode
R16624 N16623 N16624 10
D16624 N16624 0 diode
R16625 N16624 N16625 10
D16625 N16625 0 diode
R16626 N16625 N16626 10
D16626 N16626 0 diode
R16627 N16626 N16627 10
D16627 N16627 0 diode
R16628 N16627 N16628 10
D16628 N16628 0 diode
R16629 N16628 N16629 10
D16629 N16629 0 diode
R16630 N16629 N16630 10
D16630 N16630 0 diode
R16631 N16630 N16631 10
D16631 N16631 0 diode
R16632 N16631 N16632 10
D16632 N16632 0 diode
R16633 N16632 N16633 10
D16633 N16633 0 diode
R16634 N16633 N16634 10
D16634 N16634 0 diode
R16635 N16634 N16635 10
D16635 N16635 0 diode
R16636 N16635 N16636 10
D16636 N16636 0 diode
R16637 N16636 N16637 10
D16637 N16637 0 diode
R16638 N16637 N16638 10
D16638 N16638 0 diode
R16639 N16638 N16639 10
D16639 N16639 0 diode
R16640 N16639 N16640 10
D16640 N16640 0 diode
R16641 N16640 N16641 10
D16641 N16641 0 diode
R16642 N16641 N16642 10
D16642 N16642 0 diode
R16643 N16642 N16643 10
D16643 N16643 0 diode
R16644 N16643 N16644 10
D16644 N16644 0 diode
R16645 N16644 N16645 10
D16645 N16645 0 diode
R16646 N16645 N16646 10
D16646 N16646 0 diode
R16647 N16646 N16647 10
D16647 N16647 0 diode
R16648 N16647 N16648 10
D16648 N16648 0 diode
R16649 N16648 N16649 10
D16649 N16649 0 diode
R16650 N16649 N16650 10
D16650 N16650 0 diode
R16651 N16650 N16651 10
D16651 N16651 0 diode
R16652 N16651 N16652 10
D16652 N16652 0 diode
R16653 N16652 N16653 10
D16653 N16653 0 diode
R16654 N16653 N16654 10
D16654 N16654 0 diode
R16655 N16654 N16655 10
D16655 N16655 0 diode
R16656 N16655 N16656 10
D16656 N16656 0 diode
R16657 N16656 N16657 10
D16657 N16657 0 diode
R16658 N16657 N16658 10
D16658 N16658 0 diode
R16659 N16658 N16659 10
D16659 N16659 0 diode
R16660 N16659 N16660 10
D16660 N16660 0 diode
R16661 N16660 N16661 10
D16661 N16661 0 diode
R16662 N16661 N16662 10
D16662 N16662 0 diode
R16663 N16662 N16663 10
D16663 N16663 0 diode
R16664 N16663 N16664 10
D16664 N16664 0 diode
R16665 N16664 N16665 10
D16665 N16665 0 diode
R16666 N16665 N16666 10
D16666 N16666 0 diode
R16667 N16666 N16667 10
D16667 N16667 0 diode
R16668 N16667 N16668 10
D16668 N16668 0 diode
R16669 N16668 N16669 10
D16669 N16669 0 diode
R16670 N16669 N16670 10
D16670 N16670 0 diode
R16671 N16670 N16671 10
D16671 N16671 0 diode
R16672 N16671 N16672 10
D16672 N16672 0 diode
R16673 N16672 N16673 10
D16673 N16673 0 diode
R16674 N16673 N16674 10
D16674 N16674 0 diode
R16675 N16674 N16675 10
D16675 N16675 0 diode
R16676 N16675 N16676 10
D16676 N16676 0 diode
R16677 N16676 N16677 10
D16677 N16677 0 diode
R16678 N16677 N16678 10
D16678 N16678 0 diode
R16679 N16678 N16679 10
D16679 N16679 0 diode
R16680 N16679 N16680 10
D16680 N16680 0 diode
R16681 N16680 N16681 10
D16681 N16681 0 diode
R16682 N16681 N16682 10
D16682 N16682 0 diode
R16683 N16682 N16683 10
D16683 N16683 0 diode
R16684 N16683 N16684 10
D16684 N16684 0 diode
R16685 N16684 N16685 10
D16685 N16685 0 diode
R16686 N16685 N16686 10
D16686 N16686 0 diode
R16687 N16686 N16687 10
D16687 N16687 0 diode
R16688 N16687 N16688 10
D16688 N16688 0 diode
R16689 N16688 N16689 10
D16689 N16689 0 diode
R16690 N16689 N16690 10
D16690 N16690 0 diode
R16691 N16690 N16691 10
D16691 N16691 0 diode
R16692 N16691 N16692 10
D16692 N16692 0 diode
R16693 N16692 N16693 10
D16693 N16693 0 diode
R16694 N16693 N16694 10
D16694 N16694 0 diode
R16695 N16694 N16695 10
D16695 N16695 0 diode
R16696 N16695 N16696 10
D16696 N16696 0 diode
R16697 N16696 N16697 10
D16697 N16697 0 diode
R16698 N16697 N16698 10
D16698 N16698 0 diode
R16699 N16698 N16699 10
D16699 N16699 0 diode
R16700 N16699 N16700 10
D16700 N16700 0 diode
R16701 N16700 N16701 10
D16701 N16701 0 diode
R16702 N16701 N16702 10
D16702 N16702 0 diode
R16703 N16702 N16703 10
D16703 N16703 0 diode
R16704 N16703 N16704 10
D16704 N16704 0 diode
R16705 N16704 N16705 10
D16705 N16705 0 diode
R16706 N16705 N16706 10
D16706 N16706 0 diode
R16707 N16706 N16707 10
D16707 N16707 0 diode
R16708 N16707 N16708 10
D16708 N16708 0 diode
R16709 N16708 N16709 10
D16709 N16709 0 diode
R16710 N16709 N16710 10
D16710 N16710 0 diode
R16711 N16710 N16711 10
D16711 N16711 0 diode
R16712 N16711 N16712 10
D16712 N16712 0 diode
R16713 N16712 N16713 10
D16713 N16713 0 diode
R16714 N16713 N16714 10
D16714 N16714 0 diode
R16715 N16714 N16715 10
D16715 N16715 0 diode
R16716 N16715 N16716 10
D16716 N16716 0 diode
R16717 N16716 N16717 10
D16717 N16717 0 diode
R16718 N16717 N16718 10
D16718 N16718 0 diode
R16719 N16718 N16719 10
D16719 N16719 0 diode
R16720 N16719 N16720 10
D16720 N16720 0 diode
R16721 N16720 N16721 10
D16721 N16721 0 diode
R16722 N16721 N16722 10
D16722 N16722 0 diode
R16723 N16722 N16723 10
D16723 N16723 0 diode
R16724 N16723 N16724 10
D16724 N16724 0 diode
R16725 N16724 N16725 10
D16725 N16725 0 diode
R16726 N16725 N16726 10
D16726 N16726 0 diode
R16727 N16726 N16727 10
D16727 N16727 0 diode
R16728 N16727 N16728 10
D16728 N16728 0 diode
R16729 N16728 N16729 10
D16729 N16729 0 diode
R16730 N16729 N16730 10
D16730 N16730 0 diode
R16731 N16730 N16731 10
D16731 N16731 0 diode
R16732 N16731 N16732 10
D16732 N16732 0 diode
R16733 N16732 N16733 10
D16733 N16733 0 diode
R16734 N16733 N16734 10
D16734 N16734 0 diode
R16735 N16734 N16735 10
D16735 N16735 0 diode
R16736 N16735 N16736 10
D16736 N16736 0 diode
R16737 N16736 N16737 10
D16737 N16737 0 diode
R16738 N16737 N16738 10
D16738 N16738 0 diode
R16739 N16738 N16739 10
D16739 N16739 0 diode
R16740 N16739 N16740 10
D16740 N16740 0 diode
R16741 N16740 N16741 10
D16741 N16741 0 diode
R16742 N16741 N16742 10
D16742 N16742 0 diode
R16743 N16742 N16743 10
D16743 N16743 0 diode
R16744 N16743 N16744 10
D16744 N16744 0 diode
R16745 N16744 N16745 10
D16745 N16745 0 diode
R16746 N16745 N16746 10
D16746 N16746 0 diode
R16747 N16746 N16747 10
D16747 N16747 0 diode
R16748 N16747 N16748 10
D16748 N16748 0 diode
R16749 N16748 N16749 10
D16749 N16749 0 diode
R16750 N16749 N16750 10
D16750 N16750 0 diode
R16751 N16750 N16751 10
D16751 N16751 0 diode
R16752 N16751 N16752 10
D16752 N16752 0 diode
R16753 N16752 N16753 10
D16753 N16753 0 diode
R16754 N16753 N16754 10
D16754 N16754 0 diode
R16755 N16754 N16755 10
D16755 N16755 0 diode
R16756 N16755 N16756 10
D16756 N16756 0 diode
R16757 N16756 N16757 10
D16757 N16757 0 diode
R16758 N16757 N16758 10
D16758 N16758 0 diode
R16759 N16758 N16759 10
D16759 N16759 0 diode
R16760 N16759 N16760 10
D16760 N16760 0 diode
R16761 N16760 N16761 10
D16761 N16761 0 diode
R16762 N16761 N16762 10
D16762 N16762 0 diode
R16763 N16762 N16763 10
D16763 N16763 0 diode
R16764 N16763 N16764 10
D16764 N16764 0 diode
R16765 N16764 N16765 10
D16765 N16765 0 diode
R16766 N16765 N16766 10
D16766 N16766 0 diode
R16767 N16766 N16767 10
D16767 N16767 0 diode
R16768 N16767 N16768 10
D16768 N16768 0 diode
R16769 N16768 N16769 10
D16769 N16769 0 diode
R16770 N16769 N16770 10
D16770 N16770 0 diode
R16771 N16770 N16771 10
D16771 N16771 0 diode
R16772 N16771 N16772 10
D16772 N16772 0 diode
R16773 N16772 N16773 10
D16773 N16773 0 diode
R16774 N16773 N16774 10
D16774 N16774 0 diode
R16775 N16774 N16775 10
D16775 N16775 0 diode
R16776 N16775 N16776 10
D16776 N16776 0 diode
R16777 N16776 N16777 10
D16777 N16777 0 diode
R16778 N16777 N16778 10
D16778 N16778 0 diode
R16779 N16778 N16779 10
D16779 N16779 0 diode
R16780 N16779 N16780 10
D16780 N16780 0 diode
R16781 N16780 N16781 10
D16781 N16781 0 diode
R16782 N16781 N16782 10
D16782 N16782 0 diode
R16783 N16782 N16783 10
D16783 N16783 0 diode
R16784 N16783 N16784 10
D16784 N16784 0 diode
R16785 N16784 N16785 10
D16785 N16785 0 diode
R16786 N16785 N16786 10
D16786 N16786 0 diode
R16787 N16786 N16787 10
D16787 N16787 0 diode
R16788 N16787 N16788 10
D16788 N16788 0 diode
R16789 N16788 N16789 10
D16789 N16789 0 diode
R16790 N16789 N16790 10
D16790 N16790 0 diode
R16791 N16790 N16791 10
D16791 N16791 0 diode
R16792 N16791 N16792 10
D16792 N16792 0 diode
R16793 N16792 N16793 10
D16793 N16793 0 diode
R16794 N16793 N16794 10
D16794 N16794 0 diode
R16795 N16794 N16795 10
D16795 N16795 0 diode
R16796 N16795 N16796 10
D16796 N16796 0 diode
R16797 N16796 N16797 10
D16797 N16797 0 diode
R16798 N16797 N16798 10
D16798 N16798 0 diode
R16799 N16798 N16799 10
D16799 N16799 0 diode
R16800 N16799 N16800 10
D16800 N16800 0 diode
R16801 N16800 N16801 10
D16801 N16801 0 diode
R16802 N16801 N16802 10
D16802 N16802 0 diode
R16803 N16802 N16803 10
D16803 N16803 0 diode
R16804 N16803 N16804 10
D16804 N16804 0 diode
R16805 N16804 N16805 10
D16805 N16805 0 diode
R16806 N16805 N16806 10
D16806 N16806 0 diode
R16807 N16806 N16807 10
D16807 N16807 0 diode
R16808 N16807 N16808 10
D16808 N16808 0 diode
R16809 N16808 N16809 10
D16809 N16809 0 diode
R16810 N16809 N16810 10
D16810 N16810 0 diode
R16811 N16810 N16811 10
D16811 N16811 0 diode
R16812 N16811 N16812 10
D16812 N16812 0 diode
R16813 N16812 N16813 10
D16813 N16813 0 diode
R16814 N16813 N16814 10
D16814 N16814 0 diode
R16815 N16814 N16815 10
D16815 N16815 0 diode
R16816 N16815 N16816 10
D16816 N16816 0 diode
R16817 N16816 N16817 10
D16817 N16817 0 diode
R16818 N16817 N16818 10
D16818 N16818 0 diode
R16819 N16818 N16819 10
D16819 N16819 0 diode
R16820 N16819 N16820 10
D16820 N16820 0 diode
R16821 N16820 N16821 10
D16821 N16821 0 diode
R16822 N16821 N16822 10
D16822 N16822 0 diode
R16823 N16822 N16823 10
D16823 N16823 0 diode
R16824 N16823 N16824 10
D16824 N16824 0 diode
R16825 N16824 N16825 10
D16825 N16825 0 diode
R16826 N16825 N16826 10
D16826 N16826 0 diode
R16827 N16826 N16827 10
D16827 N16827 0 diode
R16828 N16827 N16828 10
D16828 N16828 0 diode
R16829 N16828 N16829 10
D16829 N16829 0 diode
R16830 N16829 N16830 10
D16830 N16830 0 diode
R16831 N16830 N16831 10
D16831 N16831 0 diode
R16832 N16831 N16832 10
D16832 N16832 0 diode
R16833 N16832 N16833 10
D16833 N16833 0 diode
R16834 N16833 N16834 10
D16834 N16834 0 diode
R16835 N16834 N16835 10
D16835 N16835 0 diode
R16836 N16835 N16836 10
D16836 N16836 0 diode
R16837 N16836 N16837 10
D16837 N16837 0 diode
R16838 N16837 N16838 10
D16838 N16838 0 diode
R16839 N16838 N16839 10
D16839 N16839 0 diode
R16840 N16839 N16840 10
D16840 N16840 0 diode
R16841 N16840 N16841 10
D16841 N16841 0 diode
R16842 N16841 N16842 10
D16842 N16842 0 diode
R16843 N16842 N16843 10
D16843 N16843 0 diode
R16844 N16843 N16844 10
D16844 N16844 0 diode
R16845 N16844 N16845 10
D16845 N16845 0 diode
R16846 N16845 N16846 10
D16846 N16846 0 diode
R16847 N16846 N16847 10
D16847 N16847 0 diode
R16848 N16847 N16848 10
D16848 N16848 0 diode
R16849 N16848 N16849 10
D16849 N16849 0 diode
R16850 N16849 N16850 10
D16850 N16850 0 diode
R16851 N16850 N16851 10
D16851 N16851 0 diode
R16852 N16851 N16852 10
D16852 N16852 0 diode
R16853 N16852 N16853 10
D16853 N16853 0 diode
R16854 N16853 N16854 10
D16854 N16854 0 diode
R16855 N16854 N16855 10
D16855 N16855 0 diode
R16856 N16855 N16856 10
D16856 N16856 0 diode
R16857 N16856 N16857 10
D16857 N16857 0 diode
R16858 N16857 N16858 10
D16858 N16858 0 diode
R16859 N16858 N16859 10
D16859 N16859 0 diode
R16860 N16859 N16860 10
D16860 N16860 0 diode
R16861 N16860 N16861 10
D16861 N16861 0 diode
R16862 N16861 N16862 10
D16862 N16862 0 diode
R16863 N16862 N16863 10
D16863 N16863 0 diode
R16864 N16863 N16864 10
D16864 N16864 0 diode
R16865 N16864 N16865 10
D16865 N16865 0 diode
R16866 N16865 N16866 10
D16866 N16866 0 diode
R16867 N16866 N16867 10
D16867 N16867 0 diode
R16868 N16867 N16868 10
D16868 N16868 0 diode
R16869 N16868 N16869 10
D16869 N16869 0 diode
R16870 N16869 N16870 10
D16870 N16870 0 diode
R16871 N16870 N16871 10
D16871 N16871 0 diode
R16872 N16871 N16872 10
D16872 N16872 0 diode
R16873 N16872 N16873 10
D16873 N16873 0 diode
R16874 N16873 N16874 10
D16874 N16874 0 diode
R16875 N16874 N16875 10
D16875 N16875 0 diode
R16876 N16875 N16876 10
D16876 N16876 0 diode
R16877 N16876 N16877 10
D16877 N16877 0 diode
R16878 N16877 N16878 10
D16878 N16878 0 diode
R16879 N16878 N16879 10
D16879 N16879 0 diode
R16880 N16879 N16880 10
D16880 N16880 0 diode
R16881 N16880 N16881 10
D16881 N16881 0 diode
R16882 N16881 N16882 10
D16882 N16882 0 diode
R16883 N16882 N16883 10
D16883 N16883 0 diode
R16884 N16883 N16884 10
D16884 N16884 0 diode
R16885 N16884 N16885 10
D16885 N16885 0 diode
R16886 N16885 N16886 10
D16886 N16886 0 diode
R16887 N16886 N16887 10
D16887 N16887 0 diode
R16888 N16887 N16888 10
D16888 N16888 0 diode
R16889 N16888 N16889 10
D16889 N16889 0 diode
R16890 N16889 N16890 10
D16890 N16890 0 diode
R16891 N16890 N16891 10
D16891 N16891 0 diode
R16892 N16891 N16892 10
D16892 N16892 0 diode
R16893 N16892 N16893 10
D16893 N16893 0 diode
R16894 N16893 N16894 10
D16894 N16894 0 diode
R16895 N16894 N16895 10
D16895 N16895 0 diode
R16896 N16895 N16896 10
D16896 N16896 0 diode
R16897 N16896 N16897 10
D16897 N16897 0 diode
R16898 N16897 N16898 10
D16898 N16898 0 diode
R16899 N16898 N16899 10
D16899 N16899 0 diode
R16900 N16899 N16900 10
D16900 N16900 0 diode
R16901 N16900 N16901 10
D16901 N16901 0 diode
R16902 N16901 N16902 10
D16902 N16902 0 diode
R16903 N16902 N16903 10
D16903 N16903 0 diode
R16904 N16903 N16904 10
D16904 N16904 0 diode
R16905 N16904 N16905 10
D16905 N16905 0 diode
R16906 N16905 N16906 10
D16906 N16906 0 diode
R16907 N16906 N16907 10
D16907 N16907 0 diode
R16908 N16907 N16908 10
D16908 N16908 0 diode
R16909 N16908 N16909 10
D16909 N16909 0 diode
R16910 N16909 N16910 10
D16910 N16910 0 diode
R16911 N16910 N16911 10
D16911 N16911 0 diode
R16912 N16911 N16912 10
D16912 N16912 0 diode
R16913 N16912 N16913 10
D16913 N16913 0 diode
R16914 N16913 N16914 10
D16914 N16914 0 diode
R16915 N16914 N16915 10
D16915 N16915 0 diode
R16916 N16915 N16916 10
D16916 N16916 0 diode
R16917 N16916 N16917 10
D16917 N16917 0 diode
R16918 N16917 N16918 10
D16918 N16918 0 diode
R16919 N16918 N16919 10
D16919 N16919 0 diode
R16920 N16919 N16920 10
D16920 N16920 0 diode
R16921 N16920 N16921 10
D16921 N16921 0 diode
R16922 N16921 N16922 10
D16922 N16922 0 diode
R16923 N16922 N16923 10
D16923 N16923 0 diode
R16924 N16923 N16924 10
D16924 N16924 0 diode
R16925 N16924 N16925 10
D16925 N16925 0 diode
R16926 N16925 N16926 10
D16926 N16926 0 diode
R16927 N16926 N16927 10
D16927 N16927 0 diode
R16928 N16927 N16928 10
D16928 N16928 0 diode
R16929 N16928 N16929 10
D16929 N16929 0 diode
R16930 N16929 N16930 10
D16930 N16930 0 diode
R16931 N16930 N16931 10
D16931 N16931 0 diode
R16932 N16931 N16932 10
D16932 N16932 0 diode
R16933 N16932 N16933 10
D16933 N16933 0 diode
R16934 N16933 N16934 10
D16934 N16934 0 diode
R16935 N16934 N16935 10
D16935 N16935 0 diode
R16936 N16935 N16936 10
D16936 N16936 0 diode
R16937 N16936 N16937 10
D16937 N16937 0 diode
R16938 N16937 N16938 10
D16938 N16938 0 diode
R16939 N16938 N16939 10
D16939 N16939 0 diode
R16940 N16939 N16940 10
D16940 N16940 0 diode
R16941 N16940 N16941 10
D16941 N16941 0 diode
R16942 N16941 N16942 10
D16942 N16942 0 diode
R16943 N16942 N16943 10
D16943 N16943 0 diode
R16944 N16943 N16944 10
D16944 N16944 0 diode
R16945 N16944 N16945 10
D16945 N16945 0 diode
R16946 N16945 N16946 10
D16946 N16946 0 diode
R16947 N16946 N16947 10
D16947 N16947 0 diode
R16948 N16947 N16948 10
D16948 N16948 0 diode
R16949 N16948 N16949 10
D16949 N16949 0 diode
R16950 N16949 N16950 10
D16950 N16950 0 diode
R16951 N16950 N16951 10
D16951 N16951 0 diode
R16952 N16951 N16952 10
D16952 N16952 0 diode
R16953 N16952 N16953 10
D16953 N16953 0 diode
R16954 N16953 N16954 10
D16954 N16954 0 diode
R16955 N16954 N16955 10
D16955 N16955 0 diode
R16956 N16955 N16956 10
D16956 N16956 0 diode
R16957 N16956 N16957 10
D16957 N16957 0 diode
R16958 N16957 N16958 10
D16958 N16958 0 diode
R16959 N16958 N16959 10
D16959 N16959 0 diode
R16960 N16959 N16960 10
D16960 N16960 0 diode
R16961 N16960 N16961 10
D16961 N16961 0 diode
R16962 N16961 N16962 10
D16962 N16962 0 diode
R16963 N16962 N16963 10
D16963 N16963 0 diode
R16964 N16963 N16964 10
D16964 N16964 0 diode
R16965 N16964 N16965 10
D16965 N16965 0 diode
R16966 N16965 N16966 10
D16966 N16966 0 diode
R16967 N16966 N16967 10
D16967 N16967 0 diode
R16968 N16967 N16968 10
D16968 N16968 0 diode
R16969 N16968 N16969 10
D16969 N16969 0 diode
R16970 N16969 N16970 10
D16970 N16970 0 diode
R16971 N16970 N16971 10
D16971 N16971 0 diode
R16972 N16971 N16972 10
D16972 N16972 0 diode
R16973 N16972 N16973 10
D16973 N16973 0 diode
R16974 N16973 N16974 10
D16974 N16974 0 diode
R16975 N16974 N16975 10
D16975 N16975 0 diode
R16976 N16975 N16976 10
D16976 N16976 0 diode
R16977 N16976 N16977 10
D16977 N16977 0 diode
R16978 N16977 N16978 10
D16978 N16978 0 diode
R16979 N16978 N16979 10
D16979 N16979 0 diode
R16980 N16979 N16980 10
D16980 N16980 0 diode
R16981 N16980 N16981 10
D16981 N16981 0 diode
R16982 N16981 N16982 10
D16982 N16982 0 diode
R16983 N16982 N16983 10
D16983 N16983 0 diode
R16984 N16983 N16984 10
D16984 N16984 0 diode
R16985 N16984 N16985 10
D16985 N16985 0 diode
R16986 N16985 N16986 10
D16986 N16986 0 diode
R16987 N16986 N16987 10
D16987 N16987 0 diode
R16988 N16987 N16988 10
D16988 N16988 0 diode
R16989 N16988 N16989 10
D16989 N16989 0 diode
R16990 N16989 N16990 10
D16990 N16990 0 diode
R16991 N16990 N16991 10
D16991 N16991 0 diode
R16992 N16991 N16992 10
D16992 N16992 0 diode
R16993 N16992 N16993 10
D16993 N16993 0 diode
R16994 N16993 N16994 10
D16994 N16994 0 diode
R16995 N16994 N16995 10
D16995 N16995 0 diode
R16996 N16995 N16996 10
D16996 N16996 0 diode
R16997 N16996 N16997 10
D16997 N16997 0 diode
R16998 N16997 N16998 10
D16998 N16998 0 diode
R16999 N16998 N16999 10
D16999 N16999 0 diode
R17000 N16999 N17000 10
D17000 N17000 0 diode
R17001 N17000 N17001 10
D17001 N17001 0 diode
R17002 N17001 N17002 10
D17002 N17002 0 diode
R17003 N17002 N17003 10
D17003 N17003 0 diode
R17004 N17003 N17004 10
D17004 N17004 0 diode
R17005 N17004 N17005 10
D17005 N17005 0 diode
R17006 N17005 N17006 10
D17006 N17006 0 diode
R17007 N17006 N17007 10
D17007 N17007 0 diode
R17008 N17007 N17008 10
D17008 N17008 0 diode
R17009 N17008 N17009 10
D17009 N17009 0 diode
R17010 N17009 N17010 10
D17010 N17010 0 diode
R17011 N17010 N17011 10
D17011 N17011 0 diode
R17012 N17011 N17012 10
D17012 N17012 0 diode
R17013 N17012 N17013 10
D17013 N17013 0 diode
R17014 N17013 N17014 10
D17014 N17014 0 diode
R17015 N17014 N17015 10
D17015 N17015 0 diode
R17016 N17015 N17016 10
D17016 N17016 0 diode
R17017 N17016 N17017 10
D17017 N17017 0 diode
R17018 N17017 N17018 10
D17018 N17018 0 diode
R17019 N17018 N17019 10
D17019 N17019 0 diode
R17020 N17019 N17020 10
D17020 N17020 0 diode
R17021 N17020 N17021 10
D17021 N17021 0 diode
R17022 N17021 N17022 10
D17022 N17022 0 diode
R17023 N17022 N17023 10
D17023 N17023 0 diode
R17024 N17023 N17024 10
D17024 N17024 0 diode
R17025 N17024 N17025 10
D17025 N17025 0 diode
R17026 N17025 N17026 10
D17026 N17026 0 diode
R17027 N17026 N17027 10
D17027 N17027 0 diode
R17028 N17027 N17028 10
D17028 N17028 0 diode
R17029 N17028 N17029 10
D17029 N17029 0 diode
R17030 N17029 N17030 10
D17030 N17030 0 diode
R17031 N17030 N17031 10
D17031 N17031 0 diode
R17032 N17031 N17032 10
D17032 N17032 0 diode
R17033 N17032 N17033 10
D17033 N17033 0 diode
R17034 N17033 N17034 10
D17034 N17034 0 diode
R17035 N17034 N17035 10
D17035 N17035 0 diode
R17036 N17035 N17036 10
D17036 N17036 0 diode
R17037 N17036 N17037 10
D17037 N17037 0 diode
R17038 N17037 N17038 10
D17038 N17038 0 diode
R17039 N17038 N17039 10
D17039 N17039 0 diode
R17040 N17039 N17040 10
D17040 N17040 0 diode
R17041 N17040 N17041 10
D17041 N17041 0 diode
R17042 N17041 N17042 10
D17042 N17042 0 diode
R17043 N17042 N17043 10
D17043 N17043 0 diode
R17044 N17043 N17044 10
D17044 N17044 0 diode
R17045 N17044 N17045 10
D17045 N17045 0 diode
R17046 N17045 N17046 10
D17046 N17046 0 diode
R17047 N17046 N17047 10
D17047 N17047 0 diode
R17048 N17047 N17048 10
D17048 N17048 0 diode
R17049 N17048 N17049 10
D17049 N17049 0 diode
R17050 N17049 N17050 10
D17050 N17050 0 diode
R17051 N17050 N17051 10
D17051 N17051 0 diode
R17052 N17051 N17052 10
D17052 N17052 0 diode
R17053 N17052 N17053 10
D17053 N17053 0 diode
R17054 N17053 N17054 10
D17054 N17054 0 diode
R17055 N17054 N17055 10
D17055 N17055 0 diode
R17056 N17055 N17056 10
D17056 N17056 0 diode
R17057 N17056 N17057 10
D17057 N17057 0 diode
R17058 N17057 N17058 10
D17058 N17058 0 diode
R17059 N17058 N17059 10
D17059 N17059 0 diode
R17060 N17059 N17060 10
D17060 N17060 0 diode
R17061 N17060 N17061 10
D17061 N17061 0 diode
R17062 N17061 N17062 10
D17062 N17062 0 diode
R17063 N17062 N17063 10
D17063 N17063 0 diode
R17064 N17063 N17064 10
D17064 N17064 0 diode
R17065 N17064 N17065 10
D17065 N17065 0 diode
R17066 N17065 N17066 10
D17066 N17066 0 diode
R17067 N17066 N17067 10
D17067 N17067 0 diode
R17068 N17067 N17068 10
D17068 N17068 0 diode
R17069 N17068 N17069 10
D17069 N17069 0 diode
R17070 N17069 N17070 10
D17070 N17070 0 diode
R17071 N17070 N17071 10
D17071 N17071 0 diode
R17072 N17071 N17072 10
D17072 N17072 0 diode
R17073 N17072 N17073 10
D17073 N17073 0 diode
R17074 N17073 N17074 10
D17074 N17074 0 diode
R17075 N17074 N17075 10
D17075 N17075 0 diode
R17076 N17075 N17076 10
D17076 N17076 0 diode
R17077 N17076 N17077 10
D17077 N17077 0 diode
R17078 N17077 N17078 10
D17078 N17078 0 diode
R17079 N17078 N17079 10
D17079 N17079 0 diode
R17080 N17079 N17080 10
D17080 N17080 0 diode
R17081 N17080 N17081 10
D17081 N17081 0 diode
R17082 N17081 N17082 10
D17082 N17082 0 diode
R17083 N17082 N17083 10
D17083 N17083 0 diode
R17084 N17083 N17084 10
D17084 N17084 0 diode
R17085 N17084 N17085 10
D17085 N17085 0 diode
R17086 N17085 N17086 10
D17086 N17086 0 diode
R17087 N17086 N17087 10
D17087 N17087 0 diode
R17088 N17087 N17088 10
D17088 N17088 0 diode
R17089 N17088 N17089 10
D17089 N17089 0 diode
R17090 N17089 N17090 10
D17090 N17090 0 diode
R17091 N17090 N17091 10
D17091 N17091 0 diode
R17092 N17091 N17092 10
D17092 N17092 0 diode
R17093 N17092 N17093 10
D17093 N17093 0 diode
R17094 N17093 N17094 10
D17094 N17094 0 diode
R17095 N17094 N17095 10
D17095 N17095 0 diode
R17096 N17095 N17096 10
D17096 N17096 0 diode
R17097 N17096 N17097 10
D17097 N17097 0 diode
R17098 N17097 N17098 10
D17098 N17098 0 diode
R17099 N17098 N17099 10
D17099 N17099 0 diode
R17100 N17099 N17100 10
D17100 N17100 0 diode
R17101 N17100 N17101 10
D17101 N17101 0 diode
R17102 N17101 N17102 10
D17102 N17102 0 diode
R17103 N17102 N17103 10
D17103 N17103 0 diode
R17104 N17103 N17104 10
D17104 N17104 0 diode
R17105 N17104 N17105 10
D17105 N17105 0 diode
R17106 N17105 N17106 10
D17106 N17106 0 diode
R17107 N17106 N17107 10
D17107 N17107 0 diode
R17108 N17107 N17108 10
D17108 N17108 0 diode
R17109 N17108 N17109 10
D17109 N17109 0 diode
R17110 N17109 N17110 10
D17110 N17110 0 diode
R17111 N17110 N17111 10
D17111 N17111 0 diode
R17112 N17111 N17112 10
D17112 N17112 0 diode
R17113 N17112 N17113 10
D17113 N17113 0 diode
R17114 N17113 N17114 10
D17114 N17114 0 diode
R17115 N17114 N17115 10
D17115 N17115 0 diode
R17116 N17115 N17116 10
D17116 N17116 0 diode
R17117 N17116 N17117 10
D17117 N17117 0 diode
R17118 N17117 N17118 10
D17118 N17118 0 diode
R17119 N17118 N17119 10
D17119 N17119 0 diode
R17120 N17119 N17120 10
D17120 N17120 0 diode
R17121 N17120 N17121 10
D17121 N17121 0 diode
R17122 N17121 N17122 10
D17122 N17122 0 diode
R17123 N17122 N17123 10
D17123 N17123 0 diode
R17124 N17123 N17124 10
D17124 N17124 0 diode
R17125 N17124 N17125 10
D17125 N17125 0 diode
R17126 N17125 N17126 10
D17126 N17126 0 diode
R17127 N17126 N17127 10
D17127 N17127 0 diode
R17128 N17127 N17128 10
D17128 N17128 0 diode
R17129 N17128 N17129 10
D17129 N17129 0 diode
R17130 N17129 N17130 10
D17130 N17130 0 diode
R17131 N17130 N17131 10
D17131 N17131 0 diode
R17132 N17131 N17132 10
D17132 N17132 0 diode
R17133 N17132 N17133 10
D17133 N17133 0 diode
R17134 N17133 N17134 10
D17134 N17134 0 diode
R17135 N17134 N17135 10
D17135 N17135 0 diode
R17136 N17135 N17136 10
D17136 N17136 0 diode
R17137 N17136 N17137 10
D17137 N17137 0 diode
R17138 N17137 N17138 10
D17138 N17138 0 diode
R17139 N17138 N17139 10
D17139 N17139 0 diode
R17140 N17139 N17140 10
D17140 N17140 0 diode
R17141 N17140 N17141 10
D17141 N17141 0 diode
R17142 N17141 N17142 10
D17142 N17142 0 diode
R17143 N17142 N17143 10
D17143 N17143 0 diode
R17144 N17143 N17144 10
D17144 N17144 0 diode
R17145 N17144 N17145 10
D17145 N17145 0 diode
R17146 N17145 N17146 10
D17146 N17146 0 diode
R17147 N17146 N17147 10
D17147 N17147 0 diode
R17148 N17147 N17148 10
D17148 N17148 0 diode
R17149 N17148 N17149 10
D17149 N17149 0 diode
R17150 N17149 N17150 10
D17150 N17150 0 diode
R17151 N17150 N17151 10
D17151 N17151 0 diode
R17152 N17151 N17152 10
D17152 N17152 0 diode
R17153 N17152 N17153 10
D17153 N17153 0 diode
R17154 N17153 N17154 10
D17154 N17154 0 diode
R17155 N17154 N17155 10
D17155 N17155 0 diode
R17156 N17155 N17156 10
D17156 N17156 0 diode
R17157 N17156 N17157 10
D17157 N17157 0 diode
R17158 N17157 N17158 10
D17158 N17158 0 diode
R17159 N17158 N17159 10
D17159 N17159 0 diode
R17160 N17159 N17160 10
D17160 N17160 0 diode
R17161 N17160 N17161 10
D17161 N17161 0 diode
R17162 N17161 N17162 10
D17162 N17162 0 diode
R17163 N17162 N17163 10
D17163 N17163 0 diode
R17164 N17163 N17164 10
D17164 N17164 0 diode
R17165 N17164 N17165 10
D17165 N17165 0 diode
R17166 N17165 N17166 10
D17166 N17166 0 diode
R17167 N17166 N17167 10
D17167 N17167 0 diode
R17168 N17167 N17168 10
D17168 N17168 0 diode
R17169 N17168 N17169 10
D17169 N17169 0 diode
R17170 N17169 N17170 10
D17170 N17170 0 diode
R17171 N17170 N17171 10
D17171 N17171 0 diode
R17172 N17171 N17172 10
D17172 N17172 0 diode
R17173 N17172 N17173 10
D17173 N17173 0 diode
R17174 N17173 N17174 10
D17174 N17174 0 diode
R17175 N17174 N17175 10
D17175 N17175 0 diode
R17176 N17175 N17176 10
D17176 N17176 0 diode
R17177 N17176 N17177 10
D17177 N17177 0 diode
R17178 N17177 N17178 10
D17178 N17178 0 diode
R17179 N17178 N17179 10
D17179 N17179 0 diode
R17180 N17179 N17180 10
D17180 N17180 0 diode
R17181 N17180 N17181 10
D17181 N17181 0 diode
R17182 N17181 N17182 10
D17182 N17182 0 diode
R17183 N17182 N17183 10
D17183 N17183 0 diode
R17184 N17183 N17184 10
D17184 N17184 0 diode
R17185 N17184 N17185 10
D17185 N17185 0 diode
R17186 N17185 N17186 10
D17186 N17186 0 diode
R17187 N17186 N17187 10
D17187 N17187 0 diode
R17188 N17187 N17188 10
D17188 N17188 0 diode
R17189 N17188 N17189 10
D17189 N17189 0 diode
R17190 N17189 N17190 10
D17190 N17190 0 diode
R17191 N17190 N17191 10
D17191 N17191 0 diode
R17192 N17191 N17192 10
D17192 N17192 0 diode
R17193 N17192 N17193 10
D17193 N17193 0 diode
R17194 N17193 N17194 10
D17194 N17194 0 diode
R17195 N17194 N17195 10
D17195 N17195 0 diode
R17196 N17195 N17196 10
D17196 N17196 0 diode
R17197 N17196 N17197 10
D17197 N17197 0 diode
R17198 N17197 N17198 10
D17198 N17198 0 diode
R17199 N17198 N17199 10
D17199 N17199 0 diode
R17200 N17199 N17200 10
D17200 N17200 0 diode
R17201 N17200 N17201 10
D17201 N17201 0 diode
R17202 N17201 N17202 10
D17202 N17202 0 diode
R17203 N17202 N17203 10
D17203 N17203 0 diode
R17204 N17203 N17204 10
D17204 N17204 0 diode
R17205 N17204 N17205 10
D17205 N17205 0 diode
R17206 N17205 N17206 10
D17206 N17206 0 diode
R17207 N17206 N17207 10
D17207 N17207 0 diode
R17208 N17207 N17208 10
D17208 N17208 0 diode
R17209 N17208 N17209 10
D17209 N17209 0 diode
R17210 N17209 N17210 10
D17210 N17210 0 diode
R17211 N17210 N17211 10
D17211 N17211 0 diode
R17212 N17211 N17212 10
D17212 N17212 0 diode
R17213 N17212 N17213 10
D17213 N17213 0 diode
R17214 N17213 N17214 10
D17214 N17214 0 diode
R17215 N17214 N17215 10
D17215 N17215 0 diode
R17216 N17215 N17216 10
D17216 N17216 0 diode
R17217 N17216 N17217 10
D17217 N17217 0 diode
R17218 N17217 N17218 10
D17218 N17218 0 diode
R17219 N17218 N17219 10
D17219 N17219 0 diode
R17220 N17219 N17220 10
D17220 N17220 0 diode
R17221 N17220 N17221 10
D17221 N17221 0 diode
R17222 N17221 N17222 10
D17222 N17222 0 diode
R17223 N17222 N17223 10
D17223 N17223 0 diode
R17224 N17223 N17224 10
D17224 N17224 0 diode
R17225 N17224 N17225 10
D17225 N17225 0 diode
R17226 N17225 N17226 10
D17226 N17226 0 diode
R17227 N17226 N17227 10
D17227 N17227 0 diode
R17228 N17227 N17228 10
D17228 N17228 0 diode
R17229 N17228 N17229 10
D17229 N17229 0 diode
R17230 N17229 N17230 10
D17230 N17230 0 diode
R17231 N17230 N17231 10
D17231 N17231 0 diode
R17232 N17231 N17232 10
D17232 N17232 0 diode
R17233 N17232 N17233 10
D17233 N17233 0 diode
R17234 N17233 N17234 10
D17234 N17234 0 diode
R17235 N17234 N17235 10
D17235 N17235 0 diode
R17236 N17235 N17236 10
D17236 N17236 0 diode
R17237 N17236 N17237 10
D17237 N17237 0 diode
R17238 N17237 N17238 10
D17238 N17238 0 diode
R17239 N17238 N17239 10
D17239 N17239 0 diode
R17240 N17239 N17240 10
D17240 N17240 0 diode
R17241 N17240 N17241 10
D17241 N17241 0 diode
R17242 N17241 N17242 10
D17242 N17242 0 diode
R17243 N17242 N17243 10
D17243 N17243 0 diode
R17244 N17243 N17244 10
D17244 N17244 0 diode
R17245 N17244 N17245 10
D17245 N17245 0 diode
R17246 N17245 N17246 10
D17246 N17246 0 diode
R17247 N17246 N17247 10
D17247 N17247 0 diode
R17248 N17247 N17248 10
D17248 N17248 0 diode
R17249 N17248 N17249 10
D17249 N17249 0 diode
R17250 N17249 N17250 10
D17250 N17250 0 diode
R17251 N17250 N17251 10
D17251 N17251 0 diode
R17252 N17251 N17252 10
D17252 N17252 0 diode
R17253 N17252 N17253 10
D17253 N17253 0 diode
R17254 N17253 N17254 10
D17254 N17254 0 diode
R17255 N17254 N17255 10
D17255 N17255 0 diode
R17256 N17255 N17256 10
D17256 N17256 0 diode
R17257 N17256 N17257 10
D17257 N17257 0 diode
R17258 N17257 N17258 10
D17258 N17258 0 diode
R17259 N17258 N17259 10
D17259 N17259 0 diode
R17260 N17259 N17260 10
D17260 N17260 0 diode
R17261 N17260 N17261 10
D17261 N17261 0 diode
R17262 N17261 N17262 10
D17262 N17262 0 diode
R17263 N17262 N17263 10
D17263 N17263 0 diode
R17264 N17263 N17264 10
D17264 N17264 0 diode
R17265 N17264 N17265 10
D17265 N17265 0 diode
R17266 N17265 N17266 10
D17266 N17266 0 diode
R17267 N17266 N17267 10
D17267 N17267 0 diode
R17268 N17267 N17268 10
D17268 N17268 0 diode
R17269 N17268 N17269 10
D17269 N17269 0 diode
R17270 N17269 N17270 10
D17270 N17270 0 diode
R17271 N17270 N17271 10
D17271 N17271 0 diode
R17272 N17271 N17272 10
D17272 N17272 0 diode
R17273 N17272 N17273 10
D17273 N17273 0 diode
R17274 N17273 N17274 10
D17274 N17274 0 diode
R17275 N17274 N17275 10
D17275 N17275 0 diode
R17276 N17275 N17276 10
D17276 N17276 0 diode
R17277 N17276 N17277 10
D17277 N17277 0 diode
R17278 N17277 N17278 10
D17278 N17278 0 diode
R17279 N17278 N17279 10
D17279 N17279 0 diode
R17280 N17279 N17280 10
D17280 N17280 0 diode
R17281 N17280 N17281 10
D17281 N17281 0 diode
R17282 N17281 N17282 10
D17282 N17282 0 diode
R17283 N17282 N17283 10
D17283 N17283 0 diode
R17284 N17283 N17284 10
D17284 N17284 0 diode
R17285 N17284 N17285 10
D17285 N17285 0 diode
R17286 N17285 N17286 10
D17286 N17286 0 diode
R17287 N17286 N17287 10
D17287 N17287 0 diode
R17288 N17287 N17288 10
D17288 N17288 0 diode
R17289 N17288 N17289 10
D17289 N17289 0 diode
R17290 N17289 N17290 10
D17290 N17290 0 diode
R17291 N17290 N17291 10
D17291 N17291 0 diode
R17292 N17291 N17292 10
D17292 N17292 0 diode
R17293 N17292 N17293 10
D17293 N17293 0 diode
R17294 N17293 N17294 10
D17294 N17294 0 diode
R17295 N17294 N17295 10
D17295 N17295 0 diode
R17296 N17295 N17296 10
D17296 N17296 0 diode
R17297 N17296 N17297 10
D17297 N17297 0 diode
R17298 N17297 N17298 10
D17298 N17298 0 diode
R17299 N17298 N17299 10
D17299 N17299 0 diode
R17300 N17299 N17300 10
D17300 N17300 0 diode
R17301 N17300 N17301 10
D17301 N17301 0 diode
R17302 N17301 N17302 10
D17302 N17302 0 diode
R17303 N17302 N17303 10
D17303 N17303 0 diode
R17304 N17303 N17304 10
D17304 N17304 0 diode
R17305 N17304 N17305 10
D17305 N17305 0 diode
R17306 N17305 N17306 10
D17306 N17306 0 diode
R17307 N17306 N17307 10
D17307 N17307 0 diode
R17308 N17307 N17308 10
D17308 N17308 0 diode
R17309 N17308 N17309 10
D17309 N17309 0 diode
R17310 N17309 N17310 10
D17310 N17310 0 diode
R17311 N17310 N17311 10
D17311 N17311 0 diode
R17312 N17311 N17312 10
D17312 N17312 0 diode
R17313 N17312 N17313 10
D17313 N17313 0 diode
R17314 N17313 N17314 10
D17314 N17314 0 diode
R17315 N17314 N17315 10
D17315 N17315 0 diode
R17316 N17315 N17316 10
D17316 N17316 0 diode
R17317 N17316 N17317 10
D17317 N17317 0 diode
R17318 N17317 N17318 10
D17318 N17318 0 diode
R17319 N17318 N17319 10
D17319 N17319 0 diode
R17320 N17319 N17320 10
D17320 N17320 0 diode
R17321 N17320 N17321 10
D17321 N17321 0 diode
R17322 N17321 N17322 10
D17322 N17322 0 diode
R17323 N17322 N17323 10
D17323 N17323 0 diode
R17324 N17323 N17324 10
D17324 N17324 0 diode
R17325 N17324 N17325 10
D17325 N17325 0 diode
R17326 N17325 N17326 10
D17326 N17326 0 diode
R17327 N17326 N17327 10
D17327 N17327 0 diode
R17328 N17327 N17328 10
D17328 N17328 0 diode
R17329 N17328 N17329 10
D17329 N17329 0 diode
R17330 N17329 N17330 10
D17330 N17330 0 diode
R17331 N17330 N17331 10
D17331 N17331 0 diode
R17332 N17331 N17332 10
D17332 N17332 0 diode
R17333 N17332 N17333 10
D17333 N17333 0 diode
R17334 N17333 N17334 10
D17334 N17334 0 diode
R17335 N17334 N17335 10
D17335 N17335 0 diode
R17336 N17335 N17336 10
D17336 N17336 0 diode
R17337 N17336 N17337 10
D17337 N17337 0 diode
R17338 N17337 N17338 10
D17338 N17338 0 diode
R17339 N17338 N17339 10
D17339 N17339 0 diode
R17340 N17339 N17340 10
D17340 N17340 0 diode
R17341 N17340 N17341 10
D17341 N17341 0 diode
R17342 N17341 N17342 10
D17342 N17342 0 diode
R17343 N17342 N17343 10
D17343 N17343 0 diode
R17344 N17343 N17344 10
D17344 N17344 0 diode
R17345 N17344 N17345 10
D17345 N17345 0 diode
R17346 N17345 N17346 10
D17346 N17346 0 diode
R17347 N17346 N17347 10
D17347 N17347 0 diode
R17348 N17347 N17348 10
D17348 N17348 0 diode
R17349 N17348 N17349 10
D17349 N17349 0 diode
R17350 N17349 N17350 10
D17350 N17350 0 diode
R17351 N17350 N17351 10
D17351 N17351 0 diode
R17352 N17351 N17352 10
D17352 N17352 0 diode
R17353 N17352 N17353 10
D17353 N17353 0 diode
R17354 N17353 N17354 10
D17354 N17354 0 diode
R17355 N17354 N17355 10
D17355 N17355 0 diode
R17356 N17355 N17356 10
D17356 N17356 0 diode
R17357 N17356 N17357 10
D17357 N17357 0 diode
R17358 N17357 N17358 10
D17358 N17358 0 diode
R17359 N17358 N17359 10
D17359 N17359 0 diode
R17360 N17359 N17360 10
D17360 N17360 0 diode
R17361 N17360 N17361 10
D17361 N17361 0 diode
R17362 N17361 N17362 10
D17362 N17362 0 diode
R17363 N17362 N17363 10
D17363 N17363 0 diode
R17364 N17363 N17364 10
D17364 N17364 0 diode
R17365 N17364 N17365 10
D17365 N17365 0 diode
R17366 N17365 N17366 10
D17366 N17366 0 diode
R17367 N17366 N17367 10
D17367 N17367 0 diode
R17368 N17367 N17368 10
D17368 N17368 0 diode
R17369 N17368 N17369 10
D17369 N17369 0 diode
R17370 N17369 N17370 10
D17370 N17370 0 diode
R17371 N17370 N17371 10
D17371 N17371 0 diode
R17372 N17371 N17372 10
D17372 N17372 0 diode
R17373 N17372 N17373 10
D17373 N17373 0 diode
R17374 N17373 N17374 10
D17374 N17374 0 diode
R17375 N17374 N17375 10
D17375 N17375 0 diode
R17376 N17375 N17376 10
D17376 N17376 0 diode
R17377 N17376 N17377 10
D17377 N17377 0 diode
R17378 N17377 N17378 10
D17378 N17378 0 diode
R17379 N17378 N17379 10
D17379 N17379 0 diode
R17380 N17379 N17380 10
D17380 N17380 0 diode
R17381 N17380 N17381 10
D17381 N17381 0 diode
R17382 N17381 N17382 10
D17382 N17382 0 diode
R17383 N17382 N17383 10
D17383 N17383 0 diode
R17384 N17383 N17384 10
D17384 N17384 0 diode
R17385 N17384 N17385 10
D17385 N17385 0 diode
R17386 N17385 N17386 10
D17386 N17386 0 diode
R17387 N17386 N17387 10
D17387 N17387 0 diode
R17388 N17387 N17388 10
D17388 N17388 0 diode
R17389 N17388 N17389 10
D17389 N17389 0 diode
R17390 N17389 N17390 10
D17390 N17390 0 diode
R17391 N17390 N17391 10
D17391 N17391 0 diode
R17392 N17391 N17392 10
D17392 N17392 0 diode
R17393 N17392 N17393 10
D17393 N17393 0 diode
R17394 N17393 N17394 10
D17394 N17394 0 diode
R17395 N17394 N17395 10
D17395 N17395 0 diode
R17396 N17395 N17396 10
D17396 N17396 0 diode
R17397 N17396 N17397 10
D17397 N17397 0 diode
R17398 N17397 N17398 10
D17398 N17398 0 diode
R17399 N17398 N17399 10
D17399 N17399 0 diode
R17400 N17399 N17400 10
D17400 N17400 0 diode
R17401 N17400 N17401 10
D17401 N17401 0 diode
R17402 N17401 N17402 10
D17402 N17402 0 diode
R17403 N17402 N17403 10
D17403 N17403 0 diode
R17404 N17403 N17404 10
D17404 N17404 0 diode
R17405 N17404 N17405 10
D17405 N17405 0 diode
R17406 N17405 N17406 10
D17406 N17406 0 diode
R17407 N17406 N17407 10
D17407 N17407 0 diode
R17408 N17407 N17408 10
D17408 N17408 0 diode
R17409 N17408 N17409 10
D17409 N17409 0 diode
R17410 N17409 N17410 10
D17410 N17410 0 diode
R17411 N17410 N17411 10
D17411 N17411 0 diode
R17412 N17411 N17412 10
D17412 N17412 0 diode
R17413 N17412 N17413 10
D17413 N17413 0 diode
R17414 N17413 N17414 10
D17414 N17414 0 diode
R17415 N17414 N17415 10
D17415 N17415 0 diode
R17416 N17415 N17416 10
D17416 N17416 0 diode
R17417 N17416 N17417 10
D17417 N17417 0 diode
R17418 N17417 N17418 10
D17418 N17418 0 diode
R17419 N17418 N17419 10
D17419 N17419 0 diode
R17420 N17419 N17420 10
D17420 N17420 0 diode
R17421 N17420 N17421 10
D17421 N17421 0 diode
R17422 N17421 N17422 10
D17422 N17422 0 diode
R17423 N17422 N17423 10
D17423 N17423 0 diode
R17424 N17423 N17424 10
D17424 N17424 0 diode
R17425 N17424 N17425 10
D17425 N17425 0 diode
R17426 N17425 N17426 10
D17426 N17426 0 diode
R17427 N17426 N17427 10
D17427 N17427 0 diode
R17428 N17427 N17428 10
D17428 N17428 0 diode
R17429 N17428 N17429 10
D17429 N17429 0 diode
R17430 N17429 N17430 10
D17430 N17430 0 diode
R17431 N17430 N17431 10
D17431 N17431 0 diode
R17432 N17431 N17432 10
D17432 N17432 0 diode
R17433 N17432 N17433 10
D17433 N17433 0 diode
R17434 N17433 N17434 10
D17434 N17434 0 diode
R17435 N17434 N17435 10
D17435 N17435 0 diode
R17436 N17435 N17436 10
D17436 N17436 0 diode
R17437 N17436 N17437 10
D17437 N17437 0 diode
R17438 N17437 N17438 10
D17438 N17438 0 diode
R17439 N17438 N17439 10
D17439 N17439 0 diode
R17440 N17439 N17440 10
D17440 N17440 0 diode
R17441 N17440 N17441 10
D17441 N17441 0 diode
R17442 N17441 N17442 10
D17442 N17442 0 diode
R17443 N17442 N17443 10
D17443 N17443 0 diode
R17444 N17443 N17444 10
D17444 N17444 0 diode
R17445 N17444 N17445 10
D17445 N17445 0 diode
R17446 N17445 N17446 10
D17446 N17446 0 diode
R17447 N17446 N17447 10
D17447 N17447 0 diode
R17448 N17447 N17448 10
D17448 N17448 0 diode
R17449 N17448 N17449 10
D17449 N17449 0 diode
R17450 N17449 N17450 10
D17450 N17450 0 diode
R17451 N17450 N17451 10
D17451 N17451 0 diode
R17452 N17451 N17452 10
D17452 N17452 0 diode
R17453 N17452 N17453 10
D17453 N17453 0 diode
R17454 N17453 N17454 10
D17454 N17454 0 diode
R17455 N17454 N17455 10
D17455 N17455 0 diode
R17456 N17455 N17456 10
D17456 N17456 0 diode
R17457 N17456 N17457 10
D17457 N17457 0 diode
R17458 N17457 N17458 10
D17458 N17458 0 diode
R17459 N17458 N17459 10
D17459 N17459 0 diode
R17460 N17459 N17460 10
D17460 N17460 0 diode
R17461 N17460 N17461 10
D17461 N17461 0 diode
R17462 N17461 N17462 10
D17462 N17462 0 diode
R17463 N17462 N17463 10
D17463 N17463 0 diode
R17464 N17463 N17464 10
D17464 N17464 0 diode
R17465 N17464 N17465 10
D17465 N17465 0 diode
R17466 N17465 N17466 10
D17466 N17466 0 diode
R17467 N17466 N17467 10
D17467 N17467 0 diode
R17468 N17467 N17468 10
D17468 N17468 0 diode
R17469 N17468 N17469 10
D17469 N17469 0 diode
R17470 N17469 N17470 10
D17470 N17470 0 diode
R17471 N17470 N17471 10
D17471 N17471 0 diode
R17472 N17471 N17472 10
D17472 N17472 0 diode
R17473 N17472 N17473 10
D17473 N17473 0 diode
R17474 N17473 N17474 10
D17474 N17474 0 diode
R17475 N17474 N17475 10
D17475 N17475 0 diode
R17476 N17475 N17476 10
D17476 N17476 0 diode
R17477 N17476 N17477 10
D17477 N17477 0 diode
R17478 N17477 N17478 10
D17478 N17478 0 diode
R17479 N17478 N17479 10
D17479 N17479 0 diode
R17480 N17479 N17480 10
D17480 N17480 0 diode
R17481 N17480 N17481 10
D17481 N17481 0 diode
R17482 N17481 N17482 10
D17482 N17482 0 diode
R17483 N17482 N17483 10
D17483 N17483 0 diode
R17484 N17483 N17484 10
D17484 N17484 0 diode
R17485 N17484 N17485 10
D17485 N17485 0 diode
R17486 N17485 N17486 10
D17486 N17486 0 diode
R17487 N17486 N17487 10
D17487 N17487 0 diode
R17488 N17487 N17488 10
D17488 N17488 0 diode
R17489 N17488 N17489 10
D17489 N17489 0 diode
R17490 N17489 N17490 10
D17490 N17490 0 diode
R17491 N17490 N17491 10
D17491 N17491 0 diode
R17492 N17491 N17492 10
D17492 N17492 0 diode
R17493 N17492 N17493 10
D17493 N17493 0 diode
R17494 N17493 N17494 10
D17494 N17494 0 diode
R17495 N17494 N17495 10
D17495 N17495 0 diode
R17496 N17495 N17496 10
D17496 N17496 0 diode
R17497 N17496 N17497 10
D17497 N17497 0 diode
R17498 N17497 N17498 10
D17498 N17498 0 diode
R17499 N17498 N17499 10
D17499 N17499 0 diode
R17500 N17499 N17500 10
D17500 N17500 0 diode
R17501 N17500 N17501 10
D17501 N17501 0 diode
R17502 N17501 N17502 10
D17502 N17502 0 diode
R17503 N17502 N17503 10
D17503 N17503 0 diode
R17504 N17503 N17504 10
D17504 N17504 0 diode
R17505 N17504 N17505 10
D17505 N17505 0 diode
R17506 N17505 N17506 10
D17506 N17506 0 diode
R17507 N17506 N17507 10
D17507 N17507 0 diode
R17508 N17507 N17508 10
D17508 N17508 0 diode
R17509 N17508 N17509 10
D17509 N17509 0 diode
R17510 N17509 N17510 10
D17510 N17510 0 diode
R17511 N17510 N17511 10
D17511 N17511 0 diode
R17512 N17511 N17512 10
D17512 N17512 0 diode
R17513 N17512 N17513 10
D17513 N17513 0 diode
R17514 N17513 N17514 10
D17514 N17514 0 diode
R17515 N17514 N17515 10
D17515 N17515 0 diode
R17516 N17515 N17516 10
D17516 N17516 0 diode
R17517 N17516 N17517 10
D17517 N17517 0 diode
R17518 N17517 N17518 10
D17518 N17518 0 diode
R17519 N17518 N17519 10
D17519 N17519 0 diode
R17520 N17519 N17520 10
D17520 N17520 0 diode
R17521 N17520 N17521 10
D17521 N17521 0 diode
R17522 N17521 N17522 10
D17522 N17522 0 diode
R17523 N17522 N17523 10
D17523 N17523 0 diode
R17524 N17523 N17524 10
D17524 N17524 0 diode
R17525 N17524 N17525 10
D17525 N17525 0 diode
R17526 N17525 N17526 10
D17526 N17526 0 diode
R17527 N17526 N17527 10
D17527 N17527 0 diode
R17528 N17527 N17528 10
D17528 N17528 0 diode
R17529 N17528 N17529 10
D17529 N17529 0 diode
R17530 N17529 N17530 10
D17530 N17530 0 diode
R17531 N17530 N17531 10
D17531 N17531 0 diode
R17532 N17531 N17532 10
D17532 N17532 0 diode
R17533 N17532 N17533 10
D17533 N17533 0 diode
R17534 N17533 N17534 10
D17534 N17534 0 diode
R17535 N17534 N17535 10
D17535 N17535 0 diode
R17536 N17535 N17536 10
D17536 N17536 0 diode
R17537 N17536 N17537 10
D17537 N17537 0 diode
R17538 N17537 N17538 10
D17538 N17538 0 diode
R17539 N17538 N17539 10
D17539 N17539 0 diode
R17540 N17539 N17540 10
D17540 N17540 0 diode
R17541 N17540 N17541 10
D17541 N17541 0 diode
R17542 N17541 N17542 10
D17542 N17542 0 diode
R17543 N17542 N17543 10
D17543 N17543 0 diode
R17544 N17543 N17544 10
D17544 N17544 0 diode
R17545 N17544 N17545 10
D17545 N17545 0 diode
R17546 N17545 N17546 10
D17546 N17546 0 diode
R17547 N17546 N17547 10
D17547 N17547 0 diode
R17548 N17547 N17548 10
D17548 N17548 0 diode
R17549 N17548 N17549 10
D17549 N17549 0 diode
R17550 N17549 N17550 10
D17550 N17550 0 diode
R17551 N17550 N17551 10
D17551 N17551 0 diode
R17552 N17551 N17552 10
D17552 N17552 0 diode
R17553 N17552 N17553 10
D17553 N17553 0 diode
R17554 N17553 N17554 10
D17554 N17554 0 diode
R17555 N17554 N17555 10
D17555 N17555 0 diode
R17556 N17555 N17556 10
D17556 N17556 0 diode
R17557 N17556 N17557 10
D17557 N17557 0 diode
R17558 N17557 N17558 10
D17558 N17558 0 diode
R17559 N17558 N17559 10
D17559 N17559 0 diode
R17560 N17559 N17560 10
D17560 N17560 0 diode
R17561 N17560 N17561 10
D17561 N17561 0 diode
R17562 N17561 N17562 10
D17562 N17562 0 diode
R17563 N17562 N17563 10
D17563 N17563 0 diode
R17564 N17563 N17564 10
D17564 N17564 0 diode
R17565 N17564 N17565 10
D17565 N17565 0 diode
R17566 N17565 N17566 10
D17566 N17566 0 diode
R17567 N17566 N17567 10
D17567 N17567 0 diode
R17568 N17567 N17568 10
D17568 N17568 0 diode
R17569 N17568 N17569 10
D17569 N17569 0 diode
R17570 N17569 N17570 10
D17570 N17570 0 diode
R17571 N17570 N17571 10
D17571 N17571 0 diode
R17572 N17571 N17572 10
D17572 N17572 0 diode
R17573 N17572 N17573 10
D17573 N17573 0 diode
R17574 N17573 N17574 10
D17574 N17574 0 diode
R17575 N17574 N17575 10
D17575 N17575 0 diode
R17576 N17575 N17576 10
D17576 N17576 0 diode
R17577 N17576 N17577 10
D17577 N17577 0 diode
R17578 N17577 N17578 10
D17578 N17578 0 diode
R17579 N17578 N17579 10
D17579 N17579 0 diode
R17580 N17579 N17580 10
D17580 N17580 0 diode
R17581 N17580 N17581 10
D17581 N17581 0 diode
R17582 N17581 N17582 10
D17582 N17582 0 diode
R17583 N17582 N17583 10
D17583 N17583 0 diode
R17584 N17583 N17584 10
D17584 N17584 0 diode
R17585 N17584 N17585 10
D17585 N17585 0 diode
R17586 N17585 N17586 10
D17586 N17586 0 diode
R17587 N17586 N17587 10
D17587 N17587 0 diode
R17588 N17587 N17588 10
D17588 N17588 0 diode
R17589 N17588 N17589 10
D17589 N17589 0 diode
R17590 N17589 N17590 10
D17590 N17590 0 diode
R17591 N17590 N17591 10
D17591 N17591 0 diode
R17592 N17591 N17592 10
D17592 N17592 0 diode
R17593 N17592 N17593 10
D17593 N17593 0 diode
R17594 N17593 N17594 10
D17594 N17594 0 diode
R17595 N17594 N17595 10
D17595 N17595 0 diode
R17596 N17595 N17596 10
D17596 N17596 0 diode
R17597 N17596 N17597 10
D17597 N17597 0 diode
R17598 N17597 N17598 10
D17598 N17598 0 diode
R17599 N17598 N17599 10
D17599 N17599 0 diode
R17600 N17599 N17600 10
D17600 N17600 0 diode
R17601 N17600 N17601 10
D17601 N17601 0 diode
R17602 N17601 N17602 10
D17602 N17602 0 diode
R17603 N17602 N17603 10
D17603 N17603 0 diode
R17604 N17603 N17604 10
D17604 N17604 0 diode
R17605 N17604 N17605 10
D17605 N17605 0 diode
R17606 N17605 N17606 10
D17606 N17606 0 diode
R17607 N17606 N17607 10
D17607 N17607 0 diode
R17608 N17607 N17608 10
D17608 N17608 0 diode
R17609 N17608 N17609 10
D17609 N17609 0 diode
R17610 N17609 N17610 10
D17610 N17610 0 diode
R17611 N17610 N17611 10
D17611 N17611 0 diode
R17612 N17611 N17612 10
D17612 N17612 0 diode
R17613 N17612 N17613 10
D17613 N17613 0 diode
R17614 N17613 N17614 10
D17614 N17614 0 diode
R17615 N17614 N17615 10
D17615 N17615 0 diode
R17616 N17615 N17616 10
D17616 N17616 0 diode
R17617 N17616 N17617 10
D17617 N17617 0 diode
R17618 N17617 N17618 10
D17618 N17618 0 diode
R17619 N17618 N17619 10
D17619 N17619 0 diode
R17620 N17619 N17620 10
D17620 N17620 0 diode
R17621 N17620 N17621 10
D17621 N17621 0 diode
R17622 N17621 N17622 10
D17622 N17622 0 diode
R17623 N17622 N17623 10
D17623 N17623 0 diode
R17624 N17623 N17624 10
D17624 N17624 0 diode
R17625 N17624 N17625 10
D17625 N17625 0 diode
R17626 N17625 N17626 10
D17626 N17626 0 diode
R17627 N17626 N17627 10
D17627 N17627 0 diode
R17628 N17627 N17628 10
D17628 N17628 0 diode
R17629 N17628 N17629 10
D17629 N17629 0 diode
R17630 N17629 N17630 10
D17630 N17630 0 diode
R17631 N17630 N17631 10
D17631 N17631 0 diode
R17632 N17631 N17632 10
D17632 N17632 0 diode
R17633 N17632 N17633 10
D17633 N17633 0 diode
R17634 N17633 N17634 10
D17634 N17634 0 diode
R17635 N17634 N17635 10
D17635 N17635 0 diode
R17636 N17635 N17636 10
D17636 N17636 0 diode
R17637 N17636 N17637 10
D17637 N17637 0 diode
R17638 N17637 N17638 10
D17638 N17638 0 diode
R17639 N17638 N17639 10
D17639 N17639 0 diode
R17640 N17639 N17640 10
D17640 N17640 0 diode
R17641 N17640 N17641 10
D17641 N17641 0 diode
R17642 N17641 N17642 10
D17642 N17642 0 diode
R17643 N17642 N17643 10
D17643 N17643 0 diode
R17644 N17643 N17644 10
D17644 N17644 0 diode
R17645 N17644 N17645 10
D17645 N17645 0 diode
R17646 N17645 N17646 10
D17646 N17646 0 diode
R17647 N17646 N17647 10
D17647 N17647 0 diode
R17648 N17647 N17648 10
D17648 N17648 0 diode
R17649 N17648 N17649 10
D17649 N17649 0 diode
R17650 N17649 N17650 10
D17650 N17650 0 diode
R17651 N17650 N17651 10
D17651 N17651 0 diode
R17652 N17651 N17652 10
D17652 N17652 0 diode
R17653 N17652 N17653 10
D17653 N17653 0 diode
R17654 N17653 N17654 10
D17654 N17654 0 diode
R17655 N17654 N17655 10
D17655 N17655 0 diode
R17656 N17655 N17656 10
D17656 N17656 0 diode
R17657 N17656 N17657 10
D17657 N17657 0 diode
R17658 N17657 N17658 10
D17658 N17658 0 diode
R17659 N17658 N17659 10
D17659 N17659 0 diode
R17660 N17659 N17660 10
D17660 N17660 0 diode
R17661 N17660 N17661 10
D17661 N17661 0 diode
R17662 N17661 N17662 10
D17662 N17662 0 diode
R17663 N17662 N17663 10
D17663 N17663 0 diode
R17664 N17663 N17664 10
D17664 N17664 0 diode
R17665 N17664 N17665 10
D17665 N17665 0 diode
R17666 N17665 N17666 10
D17666 N17666 0 diode
R17667 N17666 N17667 10
D17667 N17667 0 diode
R17668 N17667 N17668 10
D17668 N17668 0 diode
R17669 N17668 N17669 10
D17669 N17669 0 diode
R17670 N17669 N17670 10
D17670 N17670 0 diode
R17671 N17670 N17671 10
D17671 N17671 0 diode
R17672 N17671 N17672 10
D17672 N17672 0 diode
R17673 N17672 N17673 10
D17673 N17673 0 diode
R17674 N17673 N17674 10
D17674 N17674 0 diode
R17675 N17674 N17675 10
D17675 N17675 0 diode
R17676 N17675 N17676 10
D17676 N17676 0 diode
R17677 N17676 N17677 10
D17677 N17677 0 diode
R17678 N17677 N17678 10
D17678 N17678 0 diode
R17679 N17678 N17679 10
D17679 N17679 0 diode
R17680 N17679 N17680 10
D17680 N17680 0 diode
R17681 N17680 N17681 10
D17681 N17681 0 diode
R17682 N17681 N17682 10
D17682 N17682 0 diode
R17683 N17682 N17683 10
D17683 N17683 0 diode
R17684 N17683 N17684 10
D17684 N17684 0 diode
R17685 N17684 N17685 10
D17685 N17685 0 diode
R17686 N17685 N17686 10
D17686 N17686 0 diode
R17687 N17686 N17687 10
D17687 N17687 0 diode
R17688 N17687 N17688 10
D17688 N17688 0 diode
R17689 N17688 N17689 10
D17689 N17689 0 diode
R17690 N17689 N17690 10
D17690 N17690 0 diode
R17691 N17690 N17691 10
D17691 N17691 0 diode
R17692 N17691 N17692 10
D17692 N17692 0 diode
R17693 N17692 N17693 10
D17693 N17693 0 diode
R17694 N17693 N17694 10
D17694 N17694 0 diode
R17695 N17694 N17695 10
D17695 N17695 0 diode
R17696 N17695 N17696 10
D17696 N17696 0 diode
R17697 N17696 N17697 10
D17697 N17697 0 diode
R17698 N17697 N17698 10
D17698 N17698 0 diode
R17699 N17698 N17699 10
D17699 N17699 0 diode
R17700 N17699 N17700 10
D17700 N17700 0 diode
R17701 N17700 N17701 10
D17701 N17701 0 diode
R17702 N17701 N17702 10
D17702 N17702 0 diode
R17703 N17702 N17703 10
D17703 N17703 0 diode
R17704 N17703 N17704 10
D17704 N17704 0 diode
R17705 N17704 N17705 10
D17705 N17705 0 diode
R17706 N17705 N17706 10
D17706 N17706 0 diode
R17707 N17706 N17707 10
D17707 N17707 0 diode
R17708 N17707 N17708 10
D17708 N17708 0 diode
R17709 N17708 N17709 10
D17709 N17709 0 diode
R17710 N17709 N17710 10
D17710 N17710 0 diode
R17711 N17710 N17711 10
D17711 N17711 0 diode
R17712 N17711 N17712 10
D17712 N17712 0 diode
R17713 N17712 N17713 10
D17713 N17713 0 diode
R17714 N17713 N17714 10
D17714 N17714 0 diode
R17715 N17714 N17715 10
D17715 N17715 0 diode
R17716 N17715 N17716 10
D17716 N17716 0 diode
R17717 N17716 N17717 10
D17717 N17717 0 diode
R17718 N17717 N17718 10
D17718 N17718 0 diode
R17719 N17718 N17719 10
D17719 N17719 0 diode
R17720 N17719 N17720 10
D17720 N17720 0 diode
R17721 N17720 N17721 10
D17721 N17721 0 diode
R17722 N17721 N17722 10
D17722 N17722 0 diode
R17723 N17722 N17723 10
D17723 N17723 0 diode
R17724 N17723 N17724 10
D17724 N17724 0 diode
R17725 N17724 N17725 10
D17725 N17725 0 diode
R17726 N17725 N17726 10
D17726 N17726 0 diode
R17727 N17726 N17727 10
D17727 N17727 0 diode
R17728 N17727 N17728 10
D17728 N17728 0 diode
R17729 N17728 N17729 10
D17729 N17729 0 diode
R17730 N17729 N17730 10
D17730 N17730 0 diode
R17731 N17730 N17731 10
D17731 N17731 0 diode
R17732 N17731 N17732 10
D17732 N17732 0 diode
R17733 N17732 N17733 10
D17733 N17733 0 diode
R17734 N17733 N17734 10
D17734 N17734 0 diode
R17735 N17734 N17735 10
D17735 N17735 0 diode
R17736 N17735 N17736 10
D17736 N17736 0 diode
R17737 N17736 N17737 10
D17737 N17737 0 diode
R17738 N17737 N17738 10
D17738 N17738 0 diode
R17739 N17738 N17739 10
D17739 N17739 0 diode
R17740 N17739 N17740 10
D17740 N17740 0 diode
R17741 N17740 N17741 10
D17741 N17741 0 diode
R17742 N17741 N17742 10
D17742 N17742 0 diode
R17743 N17742 N17743 10
D17743 N17743 0 diode
R17744 N17743 N17744 10
D17744 N17744 0 diode
R17745 N17744 N17745 10
D17745 N17745 0 diode
R17746 N17745 N17746 10
D17746 N17746 0 diode
R17747 N17746 N17747 10
D17747 N17747 0 diode
R17748 N17747 N17748 10
D17748 N17748 0 diode
R17749 N17748 N17749 10
D17749 N17749 0 diode
R17750 N17749 N17750 10
D17750 N17750 0 diode
R17751 N17750 N17751 10
D17751 N17751 0 diode
R17752 N17751 N17752 10
D17752 N17752 0 diode
R17753 N17752 N17753 10
D17753 N17753 0 diode
R17754 N17753 N17754 10
D17754 N17754 0 diode
R17755 N17754 N17755 10
D17755 N17755 0 diode
R17756 N17755 N17756 10
D17756 N17756 0 diode
R17757 N17756 N17757 10
D17757 N17757 0 diode
R17758 N17757 N17758 10
D17758 N17758 0 diode
R17759 N17758 N17759 10
D17759 N17759 0 diode
R17760 N17759 N17760 10
D17760 N17760 0 diode
R17761 N17760 N17761 10
D17761 N17761 0 diode
R17762 N17761 N17762 10
D17762 N17762 0 diode
R17763 N17762 N17763 10
D17763 N17763 0 diode
R17764 N17763 N17764 10
D17764 N17764 0 diode
R17765 N17764 N17765 10
D17765 N17765 0 diode
R17766 N17765 N17766 10
D17766 N17766 0 diode
R17767 N17766 N17767 10
D17767 N17767 0 diode
R17768 N17767 N17768 10
D17768 N17768 0 diode
R17769 N17768 N17769 10
D17769 N17769 0 diode
R17770 N17769 N17770 10
D17770 N17770 0 diode
R17771 N17770 N17771 10
D17771 N17771 0 diode
R17772 N17771 N17772 10
D17772 N17772 0 diode
R17773 N17772 N17773 10
D17773 N17773 0 diode
R17774 N17773 N17774 10
D17774 N17774 0 diode
R17775 N17774 N17775 10
D17775 N17775 0 diode
R17776 N17775 N17776 10
D17776 N17776 0 diode
R17777 N17776 N17777 10
D17777 N17777 0 diode
R17778 N17777 N17778 10
D17778 N17778 0 diode
R17779 N17778 N17779 10
D17779 N17779 0 diode
R17780 N17779 N17780 10
D17780 N17780 0 diode
R17781 N17780 N17781 10
D17781 N17781 0 diode
R17782 N17781 N17782 10
D17782 N17782 0 diode
R17783 N17782 N17783 10
D17783 N17783 0 diode
R17784 N17783 N17784 10
D17784 N17784 0 diode
R17785 N17784 N17785 10
D17785 N17785 0 diode
R17786 N17785 N17786 10
D17786 N17786 0 diode
R17787 N17786 N17787 10
D17787 N17787 0 diode
R17788 N17787 N17788 10
D17788 N17788 0 diode
R17789 N17788 N17789 10
D17789 N17789 0 diode
R17790 N17789 N17790 10
D17790 N17790 0 diode
R17791 N17790 N17791 10
D17791 N17791 0 diode
R17792 N17791 N17792 10
D17792 N17792 0 diode
R17793 N17792 N17793 10
D17793 N17793 0 diode
R17794 N17793 N17794 10
D17794 N17794 0 diode
R17795 N17794 N17795 10
D17795 N17795 0 diode
R17796 N17795 N17796 10
D17796 N17796 0 diode
R17797 N17796 N17797 10
D17797 N17797 0 diode
R17798 N17797 N17798 10
D17798 N17798 0 diode
R17799 N17798 N17799 10
D17799 N17799 0 diode
R17800 N17799 N17800 10
D17800 N17800 0 diode
R17801 N17800 N17801 10
D17801 N17801 0 diode
R17802 N17801 N17802 10
D17802 N17802 0 diode
R17803 N17802 N17803 10
D17803 N17803 0 diode
R17804 N17803 N17804 10
D17804 N17804 0 diode
R17805 N17804 N17805 10
D17805 N17805 0 diode
R17806 N17805 N17806 10
D17806 N17806 0 diode
R17807 N17806 N17807 10
D17807 N17807 0 diode
R17808 N17807 N17808 10
D17808 N17808 0 diode
R17809 N17808 N17809 10
D17809 N17809 0 diode
R17810 N17809 N17810 10
D17810 N17810 0 diode
R17811 N17810 N17811 10
D17811 N17811 0 diode
R17812 N17811 N17812 10
D17812 N17812 0 diode
R17813 N17812 N17813 10
D17813 N17813 0 diode
R17814 N17813 N17814 10
D17814 N17814 0 diode
R17815 N17814 N17815 10
D17815 N17815 0 diode
R17816 N17815 N17816 10
D17816 N17816 0 diode
R17817 N17816 N17817 10
D17817 N17817 0 diode
R17818 N17817 N17818 10
D17818 N17818 0 diode
R17819 N17818 N17819 10
D17819 N17819 0 diode
R17820 N17819 N17820 10
D17820 N17820 0 diode
R17821 N17820 N17821 10
D17821 N17821 0 diode
R17822 N17821 N17822 10
D17822 N17822 0 diode
R17823 N17822 N17823 10
D17823 N17823 0 diode
R17824 N17823 N17824 10
D17824 N17824 0 diode
R17825 N17824 N17825 10
D17825 N17825 0 diode
R17826 N17825 N17826 10
D17826 N17826 0 diode
R17827 N17826 N17827 10
D17827 N17827 0 diode
R17828 N17827 N17828 10
D17828 N17828 0 diode
R17829 N17828 N17829 10
D17829 N17829 0 diode
R17830 N17829 N17830 10
D17830 N17830 0 diode
R17831 N17830 N17831 10
D17831 N17831 0 diode
R17832 N17831 N17832 10
D17832 N17832 0 diode
R17833 N17832 N17833 10
D17833 N17833 0 diode
R17834 N17833 N17834 10
D17834 N17834 0 diode
R17835 N17834 N17835 10
D17835 N17835 0 diode
R17836 N17835 N17836 10
D17836 N17836 0 diode
R17837 N17836 N17837 10
D17837 N17837 0 diode
R17838 N17837 N17838 10
D17838 N17838 0 diode
R17839 N17838 N17839 10
D17839 N17839 0 diode
R17840 N17839 N17840 10
D17840 N17840 0 diode
R17841 N17840 N17841 10
D17841 N17841 0 diode
R17842 N17841 N17842 10
D17842 N17842 0 diode
R17843 N17842 N17843 10
D17843 N17843 0 diode
R17844 N17843 N17844 10
D17844 N17844 0 diode
R17845 N17844 N17845 10
D17845 N17845 0 diode
R17846 N17845 N17846 10
D17846 N17846 0 diode
R17847 N17846 N17847 10
D17847 N17847 0 diode
R17848 N17847 N17848 10
D17848 N17848 0 diode
R17849 N17848 N17849 10
D17849 N17849 0 diode
R17850 N17849 N17850 10
D17850 N17850 0 diode
R17851 N17850 N17851 10
D17851 N17851 0 diode
R17852 N17851 N17852 10
D17852 N17852 0 diode
R17853 N17852 N17853 10
D17853 N17853 0 diode
R17854 N17853 N17854 10
D17854 N17854 0 diode
R17855 N17854 N17855 10
D17855 N17855 0 diode
R17856 N17855 N17856 10
D17856 N17856 0 diode
R17857 N17856 N17857 10
D17857 N17857 0 diode
R17858 N17857 N17858 10
D17858 N17858 0 diode
R17859 N17858 N17859 10
D17859 N17859 0 diode
R17860 N17859 N17860 10
D17860 N17860 0 diode
R17861 N17860 N17861 10
D17861 N17861 0 diode
R17862 N17861 N17862 10
D17862 N17862 0 diode
R17863 N17862 N17863 10
D17863 N17863 0 diode
R17864 N17863 N17864 10
D17864 N17864 0 diode
R17865 N17864 N17865 10
D17865 N17865 0 diode
R17866 N17865 N17866 10
D17866 N17866 0 diode
R17867 N17866 N17867 10
D17867 N17867 0 diode
R17868 N17867 N17868 10
D17868 N17868 0 diode
R17869 N17868 N17869 10
D17869 N17869 0 diode
R17870 N17869 N17870 10
D17870 N17870 0 diode
R17871 N17870 N17871 10
D17871 N17871 0 diode
R17872 N17871 N17872 10
D17872 N17872 0 diode
R17873 N17872 N17873 10
D17873 N17873 0 diode
R17874 N17873 N17874 10
D17874 N17874 0 diode
R17875 N17874 N17875 10
D17875 N17875 0 diode
R17876 N17875 N17876 10
D17876 N17876 0 diode
R17877 N17876 N17877 10
D17877 N17877 0 diode
R17878 N17877 N17878 10
D17878 N17878 0 diode
R17879 N17878 N17879 10
D17879 N17879 0 diode
R17880 N17879 N17880 10
D17880 N17880 0 diode
R17881 N17880 N17881 10
D17881 N17881 0 diode
R17882 N17881 N17882 10
D17882 N17882 0 diode
R17883 N17882 N17883 10
D17883 N17883 0 diode
R17884 N17883 N17884 10
D17884 N17884 0 diode
R17885 N17884 N17885 10
D17885 N17885 0 diode
R17886 N17885 N17886 10
D17886 N17886 0 diode
R17887 N17886 N17887 10
D17887 N17887 0 diode
R17888 N17887 N17888 10
D17888 N17888 0 diode
R17889 N17888 N17889 10
D17889 N17889 0 diode
R17890 N17889 N17890 10
D17890 N17890 0 diode
R17891 N17890 N17891 10
D17891 N17891 0 diode
R17892 N17891 N17892 10
D17892 N17892 0 diode
R17893 N17892 N17893 10
D17893 N17893 0 diode
R17894 N17893 N17894 10
D17894 N17894 0 diode
R17895 N17894 N17895 10
D17895 N17895 0 diode
R17896 N17895 N17896 10
D17896 N17896 0 diode
R17897 N17896 N17897 10
D17897 N17897 0 diode
R17898 N17897 N17898 10
D17898 N17898 0 diode
R17899 N17898 N17899 10
D17899 N17899 0 diode
R17900 N17899 N17900 10
D17900 N17900 0 diode
R17901 N17900 N17901 10
D17901 N17901 0 diode
R17902 N17901 N17902 10
D17902 N17902 0 diode
R17903 N17902 N17903 10
D17903 N17903 0 diode
R17904 N17903 N17904 10
D17904 N17904 0 diode
R17905 N17904 N17905 10
D17905 N17905 0 diode
R17906 N17905 N17906 10
D17906 N17906 0 diode
R17907 N17906 N17907 10
D17907 N17907 0 diode
R17908 N17907 N17908 10
D17908 N17908 0 diode
R17909 N17908 N17909 10
D17909 N17909 0 diode
R17910 N17909 N17910 10
D17910 N17910 0 diode
R17911 N17910 N17911 10
D17911 N17911 0 diode
R17912 N17911 N17912 10
D17912 N17912 0 diode
R17913 N17912 N17913 10
D17913 N17913 0 diode
R17914 N17913 N17914 10
D17914 N17914 0 diode
R17915 N17914 N17915 10
D17915 N17915 0 diode
R17916 N17915 N17916 10
D17916 N17916 0 diode
R17917 N17916 N17917 10
D17917 N17917 0 diode
R17918 N17917 N17918 10
D17918 N17918 0 diode
R17919 N17918 N17919 10
D17919 N17919 0 diode
R17920 N17919 N17920 10
D17920 N17920 0 diode
R17921 N17920 N17921 10
D17921 N17921 0 diode
R17922 N17921 N17922 10
D17922 N17922 0 diode
R17923 N17922 N17923 10
D17923 N17923 0 diode
R17924 N17923 N17924 10
D17924 N17924 0 diode
R17925 N17924 N17925 10
D17925 N17925 0 diode
R17926 N17925 N17926 10
D17926 N17926 0 diode
R17927 N17926 N17927 10
D17927 N17927 0 diode
R17928 N17927 N17928 10
D17928 N17928 0 diode
R17929 N17928 N17929 10
D17929 N17929 0 diode
R17930 N17929 N17930 10
D17930 N17930 0 diode
R17931 N17930 N17931 10
D17931 N17931 0 diode
R17932 N17931 N17932 10
D17932 N17932 0 diode
R17933 N17932 N17933 10
D17933 N17933 0 diode
R17934 N17933 N17934 10
D17934 N17934 0 diode
R17935 N17934 N17935 10
D17935 N17935 0 diode
R17936 N17935 N17936 10
D17936 N17936 0 diode
R17937 N17936 N17937 10
D17937 N17937 0 diode
R17938 N17937 N17938 10
D17938 N17938 0 diode
R17939 N17938 N17939 10
D17939 N17939 0 diode
R17940 N17939 N17940 10
D17940 N17940 0 diode
R17941 N17940 N17941 10
D17941 N17941 0 diode
R17942 N17941 N17942 10
D17942 N17942 0 diode
R17943 N17942 N17943 10
D17943 N17943 0 diode
R17944 N17943 N17944 10
D17944 N17944 0 diode
R17945 N17944 N17945 10
D17945 N17945 0 diode
R17946 N17945 N17946 10
D17946 N17946 0 diode
R17947 N17946 N17947 10
D17947 N17947 0 diode
R17948 N17947 N17948 10
D17948 N17948 0 diode
R17949 N17948 N17949 10
D17949 N17949 0 diode
R17950 N17949 N17950 10
D17950 N17950 0 diode
R17951 N17950 N17951 10
D17951 N17951 0 diode
R17952 N17951 N17952 10
D17952 N17952 0 diode
R17953 N17952 N17953 10
D17953 N17953 0 diode
R17954 N17953 N17954 10
D17954 N17954 0 diode
R17955 N17954 N17955 10
D17955 N17955 0 diode
R17956 N17955 N17956 10
D17956 N17956 0 diode
R17957 N17956 N17957 10
D17957 N17957 0 diode
R17958 N17957 N17958 10
D17958 N17958 0 diode
R17959 N17958 N17959 10
D17959 N17959 0 diode
R17960 N17959 N17960 10
D17960 N17960 0 diode
R17961 N17960 N17961 10
D17961 N17961 0 diode
R17962 N17961 N17962 10
D17962 N17962 0 diode
R17963 N17962 N17963 10
D17963 N17963 0 diode
R17964 N17963 N17964 10
D17964 N17964 0 diode
R17965 N17964 N17965 10
D17965 N17965 0 diode
R17966 N17965 N17966 10
D17966 N17966 0 diode
R17967 N17966 N17967 10
D17967 N17967 0 diode
R17968 N17967 N17968 10
D17968 N17968 0 diode
R17969 N17968 N17969 10
D17969 N17969 0 diode
R17970 N17969 N17970 10
D17970 N17970 0 diode
R17971 N17970 N17971 10
D17971 N17971 0 diode
R17972 N17971 N17972 10
D17972 N17972 0 diode
R17973 N17972 N17973 10
D17973 N17973 0 diode
R17974 N17973 N17974 10
D17974 N17974 0 diode
R17975 N17974 N17975 10
D17975 N17975 0 diode
R17976 N17975 N17976 10
D17976 N17976 0 diode
R17977 N17976 N17977 10
D17977 N17977 0 diode
R17978 N17977 N17978 10
D17978 N17978 0 diode
R17979 N17978 N17979 10
D17979 N17979 0 diode
R17980 N17979 N17980 10
D17980 N17980 0 diode
R17981 N17980 N17981 10
D17981 N17981 0 diode
R17982 N17981 N17982 10
D17982 N17982 0 diode
R17983 N17982 N17983 10
D17983 N17983 0 diode
R17984 N17983 N17984 10
D17984 N17984 0 diode
R17985 N17984 N17985 10
D17985 N17985 0 diode
R17986 N17985 N17986 10
D17986 N17986 0 diode
R17987 N17986 N17987 10
D17987 N17987 0 diode
R17988 N17987 N17988 10
D17988 N17988 0 diode
R17989 N17988 N17989 10
D17989 N17989 0 diode
R17990 N17989 N17990 10
D17990 N17990 0 diode
R17991 N17990 N17991 10
D17991 N17991 0 diode
R17992 N17991 N17992 10
D17992 N17992 0 diode
R17993 N17992 N17993 10
D17993 N17993 0 diode
R17994 N17993 N17994 10
D17994 N17994 0 diode
R17995 N17994 N17995 10
D17995 N17995 0 diode
R17996 N17995 N17996 10
D17996 N17996 0 diode
R17997 N17996 N17997 10
D17997 N17997 0 diode
R17998 N17997 N17998 10
D17998 N17998 0 diode
R17999 N17998 N17999 10
D17999 N17999 0 diode
R18000 N17999 N18000 10
D18000 N18000 0 diode
R18001 N18000 N18001 10
D18001 N18001 0 diode
R18002 N18001 N18002 10
D18002 N18002 0 diode
R18003 N18002 N18003 10
D18003 N18003 0 diode
R18004 N18003 N18004 10
D18004 N18004 0 diode
R18005 N18004 N18005 10
D18005 N18005 0 diode
R18006 N18005 N18006 10
D18006 N18006 0 diode
R18007 N18006 N18007 10
D18007 N18007 0 diode
R18008 N18007 N18008 10
D18008 N18008 0 diode
R18009 N18008 N18009 10
D18009 N18009 0 diode
R18010 N18009 N18010 10
D18010 N18010 0 diode
R18011 N18010 N18011 10
D18011 N18011 0 diode
R18012 N18011 N18012 10
D18012 N18012 0 diode
R18013 N18012 N18013 10
D18013 N18013 0 diode
R18014 N18013 N18014 10
D18014 N18014 0 diode
R18015 N18014 N18015 10
D18015 N18015 0 diode
R18016 N18015 N18016 10
D18016 N18016 0 diode
R18017 N18016 N18017 10
D18017 N18017 0 diode
R18018 N18017 N18018 10
D18018 N18018 0 diode
R18019 N18018 N18019 10
D18019 N18019 0 diode
R18020 N18019 N18020 10
D18020 N18020 0 diode
R18021 N18020 N18021 10
D18021 N18021 0 diode
R18022 N18021 N18022 10
D18022 N18022 0 diode
R18023 N18022 N18023 10
D18023 N18023 0 diode
R18024 N18023 N18024 10
D18024 N18024 0 diode
R18025 N18024 N18025 10
D18025 N18025 0 diode
R18026 N18025 N18026 10
D18026 N18026 0 diode
R18027 N18026 N18027 10
D18027 N18027 0 diode
R18028 N18027 N18028 10
D18028 N18028 0 diode
R18029 N18028 N18029 10
D18029 N18029 0 diode
R18030 N18029 N18030 10
D18030 N18030 0 diode
R18031 N18030 N18031 10
D18031 N18031 0 diode
R18032 N18031 N18032 10
D18032 N18032 0 diode
R18033 N18032 N18033 10
D18033 N18033 0 diode
R18034 N18033 N18034 10
D18034 N18034 0 diode
R18035 N18034 N18035 10
D18035 N18035 0 diode
R18036 N18035 N18036 10
D18036 N18036 0 diode
R18037 N18036 N18037 10
D18037 N18037 0 diode
R18038 N18037 N18038 10
D18038 N18038 0 diode
R18039 N18038 N18039 10
D18039 N18039 0 diode
R18040 N18039 N18040 10
D18040 N18040 0 diode
R18041 N18040 N18041 10
D18041 N18041 0 diode
R18042 N18041 N18042 10
D18042 N18042 0 diode
R18043 N18042 N18043 10
D18043 N18043 0 diode
R18044 N18043 N18044 10
D18044 N18044 0 diode
R18045 N18044 N18045 10
D18045 N18045 0 diode
R18046 N18045 N18046 10
D18046 N18046 0 diode
R18047 N18046 N18047 10
D18047 N18047 0 diode
R18048 N18047 N18048 10
D18048 N18048 0 diode
R18049 N18048 N18049 10
D18049 N18049 0 diode
R18050 N18049 N18050 10
D18050 N18050 0 diode
R18051 N18050 N18051 10
D18051 N18051 0 diode
R18052 N18051 N18052 10
D18052 N18052 0 diode
R18053 N18052 N18053 10
D18053 N18053 0 diode
R18054 N18053 N18054 10
D18054 N18054 0 diode
R18055 N18054 N18055 10
D18055 N18055 0 diode
R18056 N18055 N18056 10
D18056 N18056 0 diode
R18057 N18056 N18057 10
D18057 N18057 0 diode
R18058 N18057 N18058 10
D18058 N18058 0 diode
R18059 N18058 N18059 10
D18059 N18059 0 diode
R18060 N18059 N18060 10
D18060 N18060 0 diode
R18061 N18060 N18061 10
D18061 N18061 0 diode
R18062 N18061 N18062 10
D18062 N18062 0 diode
R18063 N18062 N18063 10
D18063 N18063 0 diode
R18064 N18063 N18064 10
D18064 N18064 0 diode
R18065 N18064 N18065 10
D18065 N18065 0 diode
R18066 N18065 N18066 10
D18066 N18066 0 diode
R18067 N18066 N18067 10
D18067 N18067 0 diode
R18068 N18067 N18068 10
D18068 N18068 0 diode
R18069 N18068 N18069 10
D18069 N18069 0 diode
R18070 N18069 N18070 10
D18070 N18070 0 diode
R18071 N18070 N18071 10
D18071 N18071 0 diode
R18072 N18071 N18072 10
D18072 N18072 0 diode
R18073 N18072 N18073 10
D18073 N18073 0 diode
R18074 N18073 N18074 10
D18074 N18074 0 diode
R18075 N18074 N18075 10
D18075 N18075 0 diode
R18076 N18075 N18076 10
D18076 N18076 0 diode
R18077 N18076 N18077 10
D18077 N18077 0 diode
R18078 N18077 N18078 10
D18078 N18078 0 diode
R18079 N18078 N18079 10
D18079 N18079 0 diode
R18080 N18079 N18080 10
D18080 N18080 0 diode
R18081 N18080 N18081 10
D18081 N18081 0 diode
R18082 N18081 N18082 10
D18082 N18082 0 diode
R18083 N18082 N18083 10
D18083 N18083 0 diode
R18084 N18083 N18084 10
D18084 N18084 0 diode
R18085 N18084 N18085 10
D18085 N18085 0 diode
R18086 N18085 N18086 10
D18086 N18086 0 diode
R18087 N18086 N18087 10
D18087 N18087 0 diode
R18088 N18087 N18088 10
D18088 N18088 0 diode
R18089 N18088 N18089 10
D18089 N18089 0 diode
R18090 N18089 N18090 10
D18090 N18090 0 diode
R18091 N18090 N18091 10
D18091 N18091 0 diode
R18092 N18091 N18092 10
D18092 N18092 0 diode
R18093 N18092 N18093 10
D18093 N18093 0 diode
R18094 N18093 N18094 10
D18094 N18094 0 diode
R18095 N18094 N18095 10
D18095 N18095 0 diode
R18096 N18095 N18096 10
D18096 N18096 0 diode
R18097 N18096 N18097 10
D18097 N18097 0 diode
R18098 N18097 N18098 10
D18098 N18098 0 diode
R18099 N18098 N18099 10
D18099 N18099 0 diode
R18100 N18099 N18100 10
D18100 N18100 0 diode
R18101 N18100 N18101 10
D18101 N18101 0 diode
R18102 N18101 N18102 10
D18102 N18102 0 diode
R18103 N18102 N18103 10
D18103 N18103 0 diode
R18104 N18103 N18104 10
D18104 N18104 0 diode
R18105 N18104 N18105 10
D18105 N18105 0 diode
R18106 N18105 N18106 10
D18106 N18106 0 diode
R18107 N18106 N18107 10
D18107 N18107 0 diode
R18108 N18107 N18108 10
D18108 N18108 0 diode
R18109 N18108 N18109 10
D18109 N18109 0 diode
R18110 N18109 N18110 10
D18110 N18110 0 diode
R18111 N18110 N18111 10
D18111 N18111 0 diode
R18112 N18111 N18112 10
D18112 N18112 0 diode
R18113 N18112 N18113 10
D18113 N18113 0 diode
R18114 N18113 N18114 10
D18114 N18114 0 diode
R18115 N18114 N18115 10
D18115 N18115 0 diode
R18116 N18115 N18116 10
D18116 N18116 0 diode
R18117 N18116 N18117 10
D18117 N18117 0 diode
R18118 N18117 N18118 10
D18118 N18118 0 diode
R18119 N18118 N18119 10
D18119 N18119 0 diode
R18120 N18119 N18120 10
D18120 N18120 0 diode
R18121 N18120 N18121 10
D18121 N18121 0 diode
R18122 N18121 N18122 10
D18122 N18122 0 diode
R18123 N18122 N18123 10
D18123 N18123 0 diode
R18124 N18123 N18124 10
D18124 N18124 0 diode
R18125 N18124 N18125 10
D18125 N18125 0 diode
R18126 N18125 N18126 10
D18126 N18126 0 diode
R18127 N18126 N18127 10
D18127 N18127 0 diode
R18128 N18127 N18128 10
D18128 N18128 0 diode
R18129 N18128 N18129 10
D18129 N18129 0 diode
R18130 N18129 N18130 10
D18130 N18130 0 diode
R18131 N18130 N18131 10
D18131 N18131 0 diode
R18132 N18131 N18132 10
D18132 N18132 0 diode
R18133 N18132 N18133 10
D18133 N18133 0 diode
R18134 N18133 N18134 10
D18134 N18134 0 diode
R18135 N18134 N18135 10
D18135 N18135 0 diode
R18136 N18135 N18136 10
D18136 N18136 0 diode
R18137 N18136 N18137 10
D18137 N18137 0 diode
R18138 N18137 N18138 10
D18138 N18138 0 diode
R18139 N18138 N18139 10
D18139 N18139 0 diode
R18140 N18139 N18140 10
D18140 N18140 0 diode
R18141 N18140 N18141 10
D18141 N18141 0 diode
R18142 N18141 N18142 10
D18142 N18142 0 diode
R18143 N18142 N18143 10
D18143 N18143 0 diode
R18144 N18143 N18144 10
D18144 N18144 0 diode
R18145 N18144 N18145 10
D18145 N18145 0 diode
R18146 N18145 N18146 10
D18146 N18146 0 diode
R18147 N18146 N18147 10
D18147 N18147 0 diode
R18148 N18147 N18148 10
D18148 N18148 0 diode
R18149 N18148 N18149 10
D18149 N18149 0 diode
R18150 N18149 N18150 10
D18150 N18150 0 diode
R18151 N18150 N18151 10
D18151 N18151 0 diode
R18152 N18151 N18152 10
D18152 N18152 0 diode
R18153 N18152 N18153 10
D18153 N18153 0 diode
R18154 N18153 N18154 10
D18154 N18154 0 diode
R18155 N18154 N18155 10
D18155 N18155 0 diode
R18156 N18155 N18156 10
D18156 N18156 0 diode
R18157 N18156 N18157 10
D18157 N18157 0 diode
R18158 N18157 N18158 10
D18158 N18158 0 diode
R18159 N18158 N18159 10
D18159 N18159 0 diode
R18160 N18159 N18160 10
D18160 N18160 0 diode
R18161 N18160 N18161 10
D18161 N18161 0 diode
R18162 N18161 N18162 10
D18162 N18162 0 diode
R18163 N18162 N18163 10
D18163 N18163 0 diode
R18164 N18163 N18164 10
D18164 N18164 0 diode
R18165 N18164 N18165 10
D18165 N18165 0 diode
R18166 N18165 N18166 10
D18166 N18166 0 diode
R18167 N18166 N18167 10
D18167 N18167 0 diode
R18168 N18167 N18168 10
D18168 N18168 0 diode
R18169 N18168 N18169 10
D18169 N18169 0 diode
R18170 N18169 N18170 10
D18170 N18170 0 diode
R18171 N18170 N18171 10
D18171 N18171 0 diode
R18172 N18171 N18172 10
D18172 N18172 0 diode
R18173 N18172 N18173 10
D18173 N18173 0 diode
R18174 N18173 N18174 10
D18174 N18174 0 diode
R18175 N18174 N18175 10
D18175 N18175 0 diode
R18176 N18175 N18176 10
D18176 N18176 0 diode
R18177 N18176 N18177 10
D18177 N18177 0 diode
R18178 N18177 N18178 10
D18178 N18178 0 diode
R18179 N18178 N18179 10
D18179 N18179 0 diode
R18180 N18179 N18180 10
D18180 N18180 0 diode
R18181 N18180 N18181 10
D18181 N18181 0 diode
R18182 N18181 N18182 10
D18182 N18182 0 diode
R18183 N18182 N18183 10
D18183 N18183 0 diode
R18184 N18183 N18184 10
D18184 N18184 0 diode
R18185 N18184 N18185 10
D18185 N18185 0 diode
R18186 N18185 N18186 10
D18186 N18186 0 diode
R18187 N18186 N18187 10
D18187 N18187 0 diode
R18188 N18187 N18188 10
D18188 N18188 0 diode
R18189 N18188 N18189 10
D18189 N18189 0 diode
R18190 N18189 N18190 10
D18190 N18190 0 diode
R18191 N18190 N18191 10
D18191 N18191 0 diode
R18192 N18191 N18192 10
D18192 N18192 0 diode
R18193 N18192 N18193 10
D18193 N18193 0 diode
R18194 N18193 N18194 10
D18194 N18194 0 diode
R18195 N18194 N18195 10
D18195 N18195 0 diode
R18196 N18195 N18196 10
D18196 N18196 0 diode
R18197 N18196 N18197 10
D18197 N18197 0 diode
R18198 N18197 N18198 10
D18198 N18198 0 diode
R18199 N18198 N18199 10
D18199 N18199 0 diode
R18200 N18199 N18200 10
D18200 N18200 0 diode
R18201 N18200 N18201 10
D18201 N18201 0 diode
R18202 N18201 N18202 10
D18202 N18202 0 diode
R18203 N18202 N18203 10
D18203 N18203 0 diode
R18204 N18203 N18204 10
D18204 N18204 0 diode
R18205 N18204 N18205 10
D18205 N18205 0 diode
R18206 N18205 N18206 10
D18206 N18206 0 diode
R18207 N18206 N18207 10
D18207 N18207 0 diode
R18208 N18207 N18208 10
D18208 N18208 0 diode
R18209 N18208 N18209 10
D18209 N18209 0 diode
R18210 N18209 N18210 10
D18210 N18210 0 diode
R18211 N18210 N18211 10
D18211 N18211 0 diode
R18212 N18211 N18212 10
D18212 N18212 0 diode
R18213 N18212 N18213 10
D18213 N18213 0 diode
R18214 N18213 N18214 10
D18214 N18214 0 diode
R18215 N18214 N18215 10
D18215 N18215 0 diode
R18216 N18215 N18216 10
D18216 N18216 0 diode
R18217 N18216 N18217 10
D18217 N18217 0 diode
R18218 N18217 N18218 10
D18218 N18218 0 diode
R18219 N18218 N18219 10
D18219 N18219 0 diode
R18220 N18219 N18220 10
D18220 N18220 0 diode
R18221 N18220 N18221 10
D18221 N18221 0 diode
R18222 N18221 N18222 10
D18222 N18222 0 diode
R18223 N18222 N18223 10
D18223 N18223 0 diode
R18224 N18223 N18224 10
D18224 N18224 0 diode
R18225 N18224 N18225 10
D18225 N18225 0 diode
R18226 N18225 N18226 10
D18226 N18226 0 diode
R18227 N18226 N18227 10
D18227 N18227 0 diode
R18228 N18227 N18228 10
D18228 N18228 0 diode
R18229 N18228 N18229 10
D18229 N18229 0 diode
R18230 N18229 N18230 10
D18230 N18230 0 diode
R18231 N18230 N18231 10
D18231 N18231 0 diode
R18232 N18231 N18232 10
D18232 N18232 0 diode
R18233 N18232 N18233 10
D18233 N18233 0 diode
R18234 N18233 N18234 10
D18234 N18234 0 diode
R18235 N18234 N18235 10
D18235 N18235 0 diode
R18236 N18235 N18236 10
D18236 N18236 0 diode
R18237 N18236 N18237 10
D18237 N18237 0 diode
R18238 N18237 N18238 10
D18238 N18238 0 diode
R18239 N18238 N18239 10
D18239 N18239 0 diode
R18240 N18239 N18240 10
D18240 N18240 0 diode
R18241 N18240 N18241 10
D18241 N18241 0 diode
R18242 N18241 N18242 10
D18242 N18242 0 diode
R18243 N18242 N18243 10
D18243 N18243 0 diode
R18244 N18243 N18244 10
D18244 N18244 0 diode
R18245 N18244 N18245 10
D18245 N18245 0 diode
R18246 N18245 N18246 10
D18246 N18246 0 diode
R18247 N18246 N18247 10
D18247 N18247 0 diode
R18248 N18247 N18248 10
D18248 N18248 0 diode
R18249 N18248 N18249 10
D18249 N18249 0 diode
R18250 N18249 N18250 10
D18250 N18250 0 diode
R18251 N18250 N18251 10
D18251 N18251 0 diode
R18252 N18251 N18252 10
D18252 N18252 0 diode
R18253 N18252 N18253 10
D18253 N18253 0 diode
R18254 N18253 N18254 10
D18254 N18254 0 diode
R18255 N18254 N18255 10
D18255 N18255 0 diode
R18256 N18255 N18256 10
D18256 N18256 0 diode
R18257 N18256 N18257 10
D18257 N18257 0 diode
R18258 N18257 N18258 10
D18258 N18258 0 diode
R18259 N18258 N18259 10
D18259 N18259 0 diode
R18260 N18259 N18260 10
D18260 N18260 0 diode
R18261 N18260 N18261 10
D18261 N18261 0 diode
R18262 N18261 N18262 10
D18262 N18262 0 diode
R18263 N18262 N18263 10
D18263 N18263 0 diode
R18264 N18263 N18264 10
D18264 N18264 0 diode
R18265 N18264 N18265 10
D18265 N18265 0 diode
R18266 N18265 N18266 10
D18266 N18266 0 diode
R18267 N18266 N18267 10
D18267 N18267 0 diode
R18268 N18267 N18268 10
D18268 N18268 0 diode
R18269 N18268 N18269 10
D18269 N18269 0 diode
R18270 N18269 N18270 10
D18270 N18270 0 diode
R18271 N18270 N18271 10
D18271 N18271 0 diode
R18272 N18271 N18272 10
D18272 N18272 0 diode
R18273 N18272 N18273 10
D18273 N18273 0 diode
R18274 N18273 N18274 10
D18274 N18274 0 diode
R18275 N18274 N18275 10
D18275 N18275 0 diode
R18276 N18275 N18276 10
D18276 N18276 0 diode
R18277 N18276 N18277 10
D18277 N18277 0 diode
R18278 N18277 N18278 10
D18278 N18278 0 diode
R18279 N18278 N18279 10
D18279 N18279 0 diode
R18280 N18279 N18280 10
D18280 N18280 0 diode
R18281 N18280 N18281 10
D18281 N18281 0 diode
R18282 N18281 N18282 10
D18282 N18282 0 diode
R18283 N18282 N18283 10
D18283 N18283 0 diode
R18284 N18283 N18284 10
D18284 N18284 0 diode
R18285 N18284 N18285 10
D18285 N18285 0 diode
R18286 N18285 N18286 10
D18286 N18286 0 diode
R18287 N18286 N18287 10
D18287 N18287 0 diode
R18288 N18287 N18288 10
D18288 N18288 0 diode
R18289 N18288 N18289 10
D18289 N18289 0 diode
R18290 N18289 N18290 10
D18290 N18290 0 diode
R18291 N18290 N18291 10
D18291 N18291 0 diode
R18292 N18291 N18292 10
D18292 N18292 0 diode
R18293 N18292 N18293 10
D18293 N18293 0 diode
R18294 N18293 N18294 10
D18294 N18294 0 diode
R18295 N18294 N18295 10
D18295 N18295 0 diode
R18296 N18295 N18296 10
D18296 N18296 0 diode
R18297 N18296 N18297 10
D18297 N18297 0 diode
R18298 N18297 N18298 10
D18298 N18298 0 diode
R18299 N18298 N18299 10
D18299 N18299 0 diode
R18300 N18299 N18300 10
D18300 N18300 0 diode
R18301 N18300 N18301 10
D18301 N18301 0 diode
R18302 N18301 N18302 10
D18302 N18302 0 diode
R18303 N18302 N18303 10
D18303 N18303 0 diode
R18304 N18303 N18304 10
D18304 N18304 0 diode
R18305 N18304 N18305 10
D18305 N18305 0 diode
R18306 N18305 N18306 10
D18306 N18306 0 diode
R18307 N18306 N18307 10
D18307 N18307 0 diode
R18308 N18307 N18308 10
D18308 N18308 0 diode
R18309 N18308 N18309 10
D18309 N18309 0 diode
R18310 N18309 N18310 10
D18310 N18310 0 diode
R18311 N18310 N18311 10
D18311 N18311 0 diode
R18312 N18311 N18312 10
D18312 N18312 0 diode
R18313 N18312 N18313 10
D18313 N18313 0 diode
R18314 N18313 N18314 10
D18314 N18314 0 diode
R18315 N18314 N18315 10
D18315 N18315 0 diode
R18316 N18315 N18316 10
D18316 N18316 0 diode
R18317 N18316 N18317 10
D18317 N18317 0 diode
R18318 N18317 N18318 10
D18318 N18318 0 diode
R18319 N18318 N18319 10
D18319 N18319 0 diode
R18320 N18319 N18320 10
D18320 N18320 0 diode
R18321 N18320 N18321 10
D18321 N18321 0 diode
R18322 N18321 N18322 10
D18322 N18322 0 diode
R18323 N18322 N18323 10
D18323 N18323 0 diode
R18324 N18323 N18324 10
D18324 N18324 0 diode
R18325 N18324 N18325 10
D18325 N18325 0 diode
R18326 N18325 N18326 10
D18326 N18326 0 diode
R18327 N18326 N18327 10
D18327 N18327 0 diode
R18328 N18327 N18328 10
D18328 N18328 0 diode
R18329 N18328 N18329 10
D18329 N18329 0 diode
R18330 N18329 N18330 10
D18330 N18330 0 diode
R18331 N18330 N18331 10
D18331 N18331 0 diode
R18332 N18331 N18332 10
D18332 N18332 0 diode
R18333 N18332 N18333 10
D18333 N18333 0 diode
R18334 N18333 N18334 10
D18334 N18334 0 diode
R18335 N18334 N18335 10
D18335 N18335 0 diode
R18336 N18335 N18336 10
D18336 N18336 0 diode
R18337 N18336 N18337 10
D18337 N18337 0 diode
R18338 N18337 N18338 10
D18338 N18338 0 diode
R18339 N18338 N18339 10
D18339 N18339 0 diode
R18340 N18339 N18340 10
D18340 N18340 0 diode
R18341 N18340 N18341 10
D18341 N18341 0 diode
R18342 N18341 N18342 10
D18342 N18342 0 diode
R18343 N18342 N18343 10
D18343 N18343 0 diode
R18344 N18343 N18344 10
D18344 N18344 0 diode
R18345 N18344 N18345 10
D18345 N18345 0 diode
R18346 N18345 N18346 10
D18346 N18346 0 diode
R18347 N18346 N18347 10
D18347 N18347 0 diode
R18348 N18347 N18348 10
D18348 N18348 0 diode
R18349 N18348 N18349 10
D18349 N18349 0 diode
R18350 N18349 N18350 10
D18350 N18350 0 diode
R18351 N18350 N18351 10
D18351 N18351 0 diode
R18352 N18351 N18352 10
D18352 N18352 0 diode
R18353 N18352 N18353 10
D18353 N18353 0 diode
R18354 N18353 N18354 10
D18354 N18354 0 diode
R18355 N18354 N18355 10
D18355 N18355 0 diode
R18356 N18355 N18356 10
D18356 N18356 0 diode
R18357 N18356 N18357 10
D18357 N18357 0 diode
R18358 N18357 N18358 10
D18358 N18358 0 diode
R18359 N18358 N18359 10
D18359 N18359 0 diode
R18360 N18359 N18360 10
D18360 N18360 0 diode
R18361 N18360 N18361 10
D18361 N18361 0 diode
R18362 N18361 N18362 10
D18362 N18362 0 diode
R18363 N18362 N18363 10
D18363 N18363 0 diode
R18364 N18363 N18364 10
D18364 N18364 0 diode
R18365 N18364 N18365 10
D18365 N18365 0 diode
R18366 N18365 N18366 10
D18366 N18366 0 diode
R18367 N18366 N18367 10
D18367 N18367 0 diode
R18368 N18367 N18368 10
D18368 N18368 0 diode
R18369 N18368 N18369 10
D18369 N18369 0 diode
R18370 N18369 N18370 10
D18370 N18370 0 diode
R18371 N18370 N18371 10
D18371 N18371 0 diode
R18372 N18371 N18372 10
D18372 N18372 0 diode
R18373 N18372 N18373 10
D18373 N18373 0 diode
R18374 N18373 N18374 10
D18374 N18374 0 diode
R18375 N18374 N18375 10
D18375 N18375 0 diode
R18376 N18375 N18376 10
D18376 N18376 0 diode
R18377 N18376 N18377 10
D18377 N18377 0 diode
R18378 N18377 N18378 10
D18378 N18378 0 diode
R18379 N18378 N18379 10
D18379 N18379 0 diode
R18380 N18379 N18380 10
D18380 N18380 0 diode
R18381 N18380 N18381 10
D18381 N18381 0 diode
R18382 N18381 N18382 10
D18382 N18382 0 diode
R18383 N18382 N18383 10
D18383 N18383 0 diode
R18384 N18383 N18384 10
D18384 N18384 0 diode
R18385 N18384 N18385 10
D18385 N18385 0 diode
R18386 N18385 N18386 10
D18386 N18386 0 diode
R18387 N18386 N18387 10
D18387 N18387 0 diode
R18388 N18387 N18388 10
D18388 N18388 0 diode
R18389 N18388 N18389 10
D18389 N18389 0 diode
R18390 N18389 N18390 10
D18390 N18390 0 diode
R18391 N18390 N18391 10
D18391 N18391 0 diode
R18392 N18391 N18392 10
D18392 N18392 0 diode
R18393 N18392 N18393 10
D18393 N18393 0 diode
R18394 N18393 N18394 10
D18394 N18394 0 diode
R18395 N18394 N18395 10
D18395 N18395 0 diode
R18396 N18395 N18396 10
D18396 N18396 0 diode
R18397 N18396 N18397 10
D18397 N18397 0 diode
R18398 N18397 N18398 10
D18398 N18398 0 diode
R18399 N18398 N18399 10
D18399 N18399 0 diode
R18400 N18399 N18400 10
D18400 N18400 0 diode
R18401 N18400 N18401 10
D18401 N18401 0 diode
R18402 N18401 N18402 10
D18402 N18402 0 diode
R18403 N18402 N18403 10
D18403 N18403 0 diode
R18404 N18403 N18404 10
D18404 N18404 0 diode
R18405 N18404 N18405 10
D18405 N18405 0 diode
R18406 N18405 N18406 10
D18406 N18406 0 diode
R18407 N18406 N18407 10
D18407 N18407 0 diode
R18408 N18407 N18408 10
D18408 N18408 0 diode
R18409 N18408 N18409 10
D18409 N18409 0 diode
R18410 N18409 N18410 10
D18410 N18410 0 diode
R18411 N18410 N18411 10
D18411 N18411 0 diode
R18412 N18411 N18412 10
D18412 N18412 0 diode
R18413 N18412 N18413 10
D18413 N18413 0 diode
R18414 N18413 N18414 10
D18414 N18414 0 diode
R18415 N18414 N18415 10
D18415 N18415 0 diode
R18416 N18415 N18416 10
D18416 N18416 0 diode
R18417 N18416 N18417 10
D18417 N18417 0 diode
R18418 N18417 N18418 10
D18418 N18418 0 diode
R18419 N18418 N18419 10
D18419 N18419 0 diode
R18420 N18419 N18420 10
D18420 N18420 0 diode
R18421 N18420 N18421 10
D18421 N18421 0 diode
R18422 N18421 N18422 10
D18422 N18422 0 diode
R18423 N18422 N18423 10
D18423 N18423 0 diode
R18424 N18423 N18424 10
D18424 N18424 0 diode
R18425 N18424 N18425 10
D18425 N18425 0 diode
R18426 N18425 N18426 10
D18426 N18426 0 diode
R18427 N18426 N18427 10
D18427 N18427 0 diode
R18428 N18427 N18428 10
D18428 N18428 0 diode
R18429 N18428 N18429 10
D18429 N18429 0 diode
R18430 N18429 N18430 10
D18430 N18430 0 diode
R18431 N18430 N18431 10
D18431 N18431 0 diode
R18432 N18431 N18432 10
D18432 N18432 0 diode
R18433 N18432 N18433 10
D18433 N18433 0 diode
R18434 N18433 N18434 10
D18434 N18434 0 diode
R18435 N18434 N18435 10
D18435 N18435 0 diode
R18436 N18435 N18436 10
D18436 N18436 0 diode
R18437 N18436 N18437 10
D18437 N18437 0 diode
R18438 N18437 N18438 10
D18438 N18438 0 diode
R18439 N18438 N18439 10
D18439 N18439 0 diode
R18440 N18439 N18440 10
D18440 N18440 0 diode
R18441 N18440 N18441 10
D18441 N18441 0 diode
R18442 N18441 N18442 10
D18442 N18442 0 diode
R18443 N18442 N18443 10
D18443 N18443 0 diode
R18444 N18443 N18444 10
D18444 N18444 0 diode
R18445 N18444 N18445 10
D18445 N18445 0 diode
R18446 N18445 N18446 10
D18446 N18446 0 diode
R18447 N18446 N18447 10
D18447 N18447 0 diode
R18448 N18447 N18448 10
D18448 N18448 0 diode
R18449 N18448 N18449 10
D18449 N18449 0 diode
R18450 N18449 N18450 10
D18450 N18450 0 diode
R18451 N18450 N18451 10
D18451 N18451 0 diode
R18452 N18451 N18452 10
D18452 N18452 0 diode
R18453 N18452 N18453 10
D18453 N18453 0 diode
R18454 N18453 N18454 10
D18454 N18454 0 diode
R18455 N18454 N18455 10
D18455 N18455 0 diode
R18456 N18455 N18456 10
D18456 N18456 0 diode
R18457 N18456 N18457 10
D18457 N18457 0 diode
R18458 N18457 N18458 10
D18458 N18458 0 diode
R18459 N18458 N18459 10
D18459 N18459 0 diode
R18460 N18459 N18460 10
D18460 N18460 0 diode
R18461 N18460 N18461 10
D18461 N18461 0 diode
R18462 N18461 N18462 10
D18462 N18462 0 diode
R18463 N18462 N18463 10
D18463 N18463 0 diode
R18464 N18463 N18464 10
D18464 N18464 0 diode
R18465 N18464 N18465 10
D18465 N18465 0 diode
R18466 N18465 N18466 10
D18466 N18466 0 diode
R18467 N18466 N18467 10
D18467 N18467 0 diode
R18468 N18467 N18468 10
D18468 N18468 0 diode
R18469 N18468 N18469 10
D18469 N18469 0 diode
R18470 N18469 N18470 10
D18470 N18470 0 diode
R18471 N18470 N18471 10
D18471 N18471 0 diode
R18472 N18471 N18472 10
D18472 N18472 0 diode
R18473 N18472 N18473 10
D18473 N18473 0 diode
R18474 N18473 N18474 10
D18474 N18474 0 diode
R18475 N18474 N18475 10
D18475 N18475 0 diode
R18476 N18475 N18476 10
D18476 N18476 0 diode
R18477 N18476 N18477 10
D18477 N18477 0 diode
R18478 N18477 N18478 10
D18478 N18478 0 diode
R18479 N18478 N18479 10
D18479 N18479 0 diode
R18480 N18479 N18480 10
D18480 N18480 0 diode
R18481 N18480 N18481 10
D18481 N18481 0 diode
R18482 N18481 N18482 10
D18482 N18482 0 diode
R18483 N18482 N18483 10
D18483 N18483 0 diode
R18484 N18483 N18484 10
D18484 N18484 0 diode
R18485 N18484 N18485 10
D18485 N18485 0 diode
R18486 N18485 N18486 10
D18486 N18486 0 diode
R18487 N18486 N18487 10
D18487 N18487 0 diode
R18488 N18487 N18488 10
D18488 N18488 0 diode
R18489 N18488 N18489 10
D18489 N18489 0 diode
R18490 N18489 N18490 10
D18490 N18490 0 diode
R18491 N18490 N18491 10
D18491 N18491 0 diode
R18492 N18491 N18492 10
D18492 N18492 0 diode
R18493 N18492 N18493 10
D18493 N18493 0 diode
R18494 N18493 N18494 10
D18494 N18494 0 diode
R18495 N18494 N18495 10
D18495 N18495 0 diode
R18496 N18495 N18496 10
D18496 N18496 0 diode
R18497 N18496 N18497 10
D18497 N18497 0 diode
R18498 N18497 N18498 10
D18498 N18498 0 diode
R18499 N18498 N18499 10
D18499 N18499 0 diode
R18500 N18499 N18500 10
D18500 N18500 0 diode
R18501 N18500 N18501 10
D18501 N18501 0 diode
R18502 N18501 N18502 10
D18502 N18502 0 diode
R18503 N18502 N18503 10
D18503 N18503 0 diode
R18504 N18503 N18504 10
D18504 N18504 0 diode
R18505 N18504 N18505 10
D18505 N18505 0 diode
R18506 N18505 N18506 10
D18506 N18506 0 diode
R18507 N18506 N18507 10
D18507 N18507 0 diode
R18508 N18507 N18508 10
D18508 N18508 0 diode
R18509 N18508 N18509 10
D18509 N18509 0 diode
R18510 N18509 N18510 10
D18510 N18510 0 diode
R18511 N18510 N18511 10
D18511 N18511 0 diode
R18512 N18511 N18512 10
D18512 N18512 0 diode
R18513 N18512 N18513 10
D18513 N18513 0 diode
R18514 N18513 N18514 10
D18514 N18514 0 diode
R18515 N18514 N18515 10
D18515 N18515 0 diode
R18516 N18515 N18516 10
D18516 N18516 0 diode
R18517 N18516 N18517 10
D18517 N18517 0 diode
R18518 N18517 N18518 10
D18518 N18518 0 diode
R18519 N18518 N18519 10
D18519 N18519 0 diode
R18520 N18519 N18520 10
D18520 N18520 0 diode
R18521 N18520 N18521 10
D18521 N18521 0 diode
R18522 N18521 N18522 10
D18522 N18522 0 diode
R18523 N18522 N18523 10
D18523 N18523 0 diode
R18524 N18523 N18524 10
D18524 N18524 0 diode
R18525 N18524 N18525 10
D18525 N18525 0 diode
R18526 N18525 N18526 10
D18526 N18526 0 diode
R18527 N18526 N18527 10
D18527 N18527 0 diode
R18528 N18527 N18528 10
D18528 N18528 0 diode
R18529 N18528 N18529 10
D18529 N18529 0 diode
R18530 N18529 N18530 10
D18530 N18530 0 diode
R18531 N18530 N18531 10
D18531 N18531 0 diode
R18532 N18531 N18532 10
D18532 N18532 0 diode
R18533 N18532 N18533 10
D18533 N18533 0 diode
R18534 N18533 N18534 10
D18534 N18534 0 diode
R18535 N18534 N18535 10
D18535 N18535 0 diode
R18536 N18535 N18536 10
D18536 N18536 0 diode
R18537 N18536 N18537 10
D18537 N18537 0 diode
R18538 N18537 N18538 10
D18538 N18538 0 diode
R18539 N18538 N18539 10
D18539 N18539 0 diode
R18540 N18539 N18540 10
D18540 N18540 0 diode
R18541 N18540 N18541 10
D18541 N18541 0 diode
R18542 N18541 N18542 10
D18542 N18542 0 diode
R18543 N18542 N18543 10
D18543 N18543 0 diode
R18544 N18543 N18544 10
D18544 N18544 0 diode
R18545 N18544 N18545 10
D18545 N18545 0 diode
R18546 N18545 N18546 10
D18546 N18546 0 diode
R18547 N18546 N18547 10
D18547 N18547 0 diode
R18548 N18547 N18548 10
D18548 N18548 0 diode
R18549 N18548 N18549 10
D18549 N18549 0 diode
R18550 N18549 N18550 10
D18550 N18550 0 diode
R18551 N18550 N18551 10
D18551 N18551 0 diode
R18552 N18551 N18552 10
D18552 N18552 0 diode
R18553 N18552 N18553 10
D18553 N18553 0 diode
R18554 N18553 N18554 10
D18554 N18554 0 diode
R18555 N18554 N18555 10
D18555 N18555 0 diode
R18556 N18555 N18556 10
D18556 N18556 0 diode
R18557 N18556 N18557 10
D18557 N18557 0 diode
R18558 N18557 N18558 10
D18558 N18558 0 diode
R18559 N18558 N18559 10
D18559 N18559 0 diode
R18560 N18559 N18560 10
D18560 N18560 0 diode
R18561 N18560 N18561 10
D18561 N18561 0 diode
R18562 N18561 N18562 10
D18562 N18562 0 diode
R18563 N18562 N18563 10
D18563 N18563 0 diode
R18564 N18563 N18564 10
D18564 N18564 0 diode
R18565 N18564 N18565 10
D18565 N18565 0 diode
R18566 N18565 N18566 10
D18566 N18566 0 diode
R18567 N18566 N18567 10
D18567 N18567 0 diode
R18568 N18567 N18568 10
D18568 N18568 0 diode
R18569 N18568 N18569 10
D18569 N18569 0 diode
R18570 N18569 N18570 10
D18570 N18570 0 diode
R18571 N18570 N18571 10
D18571 N18571 0 diode
R18572 N18571 N18572 10
D18572 N18572 0 diode
R18573 N18572 N18573 10
D18573 N18573 0 diode
R18574 N18573 N18574 10
D18574 N18574 0 diode
R18575 N18574 N18575 10
D18575 N18575 0 diode
R18576 N18575 N18576 10
D18576 N18576 0 diode
R18577 N18576 N18577 10
D18577 N18577 0 diode
R18578 N18577 N18578 10
D18578 N18578 0 diode
R18579 N18578 N18579 10
D18579 N18579 0 diode
R18580 N18579 N18580 10
D18580 N18580 0 diode
R18581 N18580 N18581 10
D18581 N18581 0 diode
R18582 N18581 N18582 10
D18582 N18582 0 diode
R18583 N18582 N18583 10
D18583 N18583 0 diode
R18584 N18583 N18584 10
D18584 N18584 0 diode
R18585 N18584 N18585 10
D18585 N18585 0 diode
R18586 N18585 N18586 10
D18586 N18586 0 diode
R18587 N18586 N18587 10
D18587 N18587 0 diode
R18588 N18587 N18588 10
D18588 N18588 0 diode
R18589 N18588 N18589 10
D18589 N18589 0 diode
R18590 N18589 N18590 10
D18590 N18590 0 diode
R18591 N18590 N18591 10
D18591 N18591 0 diode
R18592 N18591 N18592 10
D18592 N18592 0 diode
R18593 N18592 N18593 10
D18593 N18593 0 diode
R18594 N18593 N18594 10
D18594 N18594 0 diode
R18595 N18594 N18595 10
D18595 N18595 0 diode
R18596 N18595 N18596 10
D18596 N18596 0 diode
R18597 N18596 N18597 10
D18597 N18597 0 diode
R18598 N18597 N18598 10
D18598 N18598 0 diode
R18599 N18598 N18599 10
D18599 N18599 0 diode
R18600 N18599 N18600 10
D18600 N18600 0 diode
R18601 N18600 N18601 10
D18601 N18601 0 diode
R18602 N18601 N18602 10
D18602 N18602 0 diode
R18603 N18602 N18603 10
D18603 N18603 0 diode
R18604 N18603 N18604 10
D18604 N18604 0 diode
R18605 N18604 N18605 10
D18605 N18605 0 diode
R18606 N18605 N18606 10
D18606 N18606 0 diode
R18607 N18606 N18607 10
D18607 N18607 0 diode
R18608 N18607 N18608 10
D18608 N18608 0 diode
R18609 N18608 N18609 10
D18609 N18609 0 diode
R18610 N18609 N18610 10
D18610 N18610 0 diode
R18611 N18610 N18611 10
D18611 N18611 0 diode
R18612 N18611 N18612 10
D18612 N18612 0 diode
R18613 N18612 N18613 10
D18613 N18613 0 diode
R18614 N18613 N18614 10
D18614 N18614 0 diode
R18615 N18614 N18615 10
D18615 N18615 0 diode
R18616 N18615 N18616 10
D18616 N18616 0 diode
R18617 N18616 N18617 10
D18617 N18617 0 diode
R18618 N18617 N18618 10
D18618 N18618 0 diode
R18619 N18618 N18619 10
D18619 N18619 0 diode
R18620 N18619 N18620 10
D18620 N18620 0 diode
R18621 N18620 N18621 10
D18621 N18621 0 diode
R18622 N18621 N18622 10
D18622 N18622 0 diode
R18623 N18622 N18623 10
D18623 N18623 0 diode
R18624 N18623 N18624 10
D18624 N18624 0 diode
R18625 N18624 N18625 10
D18625 N18625 0 diode
R18626 N18625 N18626 10
D18626 N18626 0 diode
R18627 N18626 N18627 10
D18627 N18627 0 diode
R18628 N18627 N18628 10
D18628 N18628 0 diode
R18629 N18628 N18629 10
D18629 N18629 0 diode
R18630 N18629 N18630 10
D18630 N18630 0 diode
R18631 N18630 N18631 10
D18631 N18631 0 diode
R18632 N18631 N18632 10
D18632 N18632 0 diode
R18633 N18632 N18633 10
D18633 N18633 0 diode
R18634 N18633 N18634 10
D18634 N18634 0 diode
R18635 N18634 N18635 10
D18635 N18635 0 diode
R18636 N18635 N18636 10
D18636 N18636 0 diode
R18637 N18636 N18637 10
D18637 N18637 0 diode
R18638 N18637 N18638 10
D18638 N18638 0 diode
R18639 N18638 N18639 10
D18639 N18639 0 diode
R18640 N18639 N18640 10
D18640 N18640 0 diode
R18641 N18640 N18641 10
D18641 N18641 0 diode
R18642 N18641 N18642 10
D18642 N18642 0 diode
R18643 N18642 N18643 10
D18643 N18643 0 diode
R18644 N18643 N18644 10
D18644 N18644 0 diode
R18645 N18644 N18645 10
D18645 N18645 0 diode
R18646 N18645 N18646 10
D18646 N18646 0 diode
R18647 N18646 N18647 10
D18647 N18647 0 diode
R18648 N18647 N18648 10
D18648 N18648 0 diode
R18649 N18648 N18649 10
D18649 N18649 0 diode
R18650 N18649 N18650 10
D18650 N18650 0 diode
R18651 N18650 N18651 10
D18651 N18651 0 diode
R18652 N18651 N18652 10
D18652 N18652 0 diode
R18653 N18652 N18653 10
D18653 N18653 0 diode
R18654 N18653 N18654 10
D18654 N18654 0 diode
R18655 N18654 N18655 10
D18655 N18655 0 diode
R18656 N18655 N18656 10
D18656 N18656 0 diode
R18657 N18656 N18657 10
D18657 N18657 0 diode
R18658 N18657 N18658 10
D18658 N18658 0 diode
R18659 N18658 N18659 10
D18659 N18659 0 diode
R18660 N18659 N18660 10
D18660 N18660 0 diode
R18661 N18660 N18661 10
D18661 N18661 0 diode
R18662 N18661 N18662 10
D18662 N18662 0 diode
R18663 N18662 N18663 10
D18663 N18663 0 diode
R18664 N18663 N18664 10
D18664 N18664 0 diode
R18665 N18664 N18665 10
D18665 N18665 0 diode
R18666 N18665 N18666 10
D18666 N18666 0 diode
R18667 N18666 N18667 10
D18667 N18667 0 diode
R18668 N18667 N18668 10
D18668 N18668 0 diode
R18669 N18668 N18669 10
D18669 N18669 0 diode
R18670 N18669 N18670 10
D18670 N18670 0 diode
R18671 N18670 N18671 10
D18671 N18671 0 diode
R18672 N18671 N18672 10
D18672 N18672 0 diode
R18673 N18672 N18673 10
D18673 N18673 0 diode
R18674 N18673 N18674 10
D18674 N18674 0 diode
R18675 N18674 N18675 10
D18675 N18675 0 diode
R18676 N18675 N18676 10
D18676 N18676 0 diode
R18677 N18676 N18677 10
D18677 N18677 0 diode
R18678 N18677 N18678 10
D18678 N18678 0 diode
R18679 N18678 N18679 10
D18679 N18679 0 diode
R18680 N18679 N18680 10
D18680 N18680 0 diode
R18681 N18680 N18681 10
D18681 N18681 0 diode
R18682 N18681 N18682 10
D18682 N18682 0 diode
R18683 N18682 N18683 10
D18683 N18683 0 diode
R18684 N18683 N18684 10
D18684 N18684 0 diode
R18685 N18684 N18685 10
D18685 N18685 0 diode
R18686 N18685 N18686 10
D18686 N18686 0 diode
R18687 N18686 N18687 10
D18687 N18687 0 diode
R18688 N18687 N18688 10
D18688 N18688 0 diode
R18689 N18688 N18689 10
D18689 N18689 0 diode
R18690 N18689 N18690 10
D18690 N18690 0 diode
R18691 N18690 N18691 10
D18691 N18691 0 diode
R18692 N18691 N18692 10
D18692 N18692 0 diode
R18693 N18692 N18693 10
D18693 N18693 0 diode
R18694 N18693 N18694 10
D18694 N18694 0 diode
R18695 N18694 N18695 10
D18695 N18695 0 diode
R18696 N18695 N18696 10
D18696 N18696 0 diode
R18697 N18696 N18697 10
D18697 N18697 0 diode
R18698 N18697 N18698 10
D18698 N18698 0 diode
R18699 N18698 N18699 10
D18699 N18699 0 diode
R18700 N18699 N18700 10
D18700 N18700 0 diode
R18701 N18700 N18701 10
D18701 N18701 0 diode
R18702 N18701 N18702 10
D18702 N18702 0 diode
R18703 N18702 N18703 10
D18703 N18703 0 diode
R18704 N18703 N18704 10
D18704 N18704 0 diode
R18705 N18704 N18705 10
D18705 N18705 0 diode
R18706 N18705 N18706 10
D18706 N18706 0 diode
R18707 N18706 N18707 10
D18707 N18707 0 diode
R18708 N18707 N18708 10
D18708 N18708 0 diode
R18709 N18708 N18709 10
D18709 N18709 0 diode
R18710 N18709 N18710 10
D18710 N18710 0 diode
R18711 N18710 N18711 10
D18711 N18711 0 diode
R18712 N18711 N18712 10
D18712 N18712 0 diode
R18713 N18712 N18713 10
D18713 N18713 0 diode
R18714 N18713 N18714 10
D18714 N18714 0 diode
R18715 N18714 N18715 10
D18715 N18715 0 diode
R18716 N18715 N18716 10
D18716 N18716 0 diode
R18717 N18716 N18717 10
D18717 N18717 0 diode
R18718 N18717 N18718 10
D18718 N18718 0 diode
R18719 N18718 N18719 10
D18719 N18719 0 diode
R18720 N18719 N18720 10
D18720 N18720 0 diode
R18721 N18720 N18721 10
D18721 N18721 0 diode
R18722 N18721 N18722 10
D18722 N18722 0 diode
R18723 N18722 N18723 10
D18723 N18723 0 diode
R18724 N18723 N18724 10
D18724 N18724 0 diode
R18725 N18724 N18725 10
D18725 N18725 0 diode
R18726 N18725 N18726 10
D18726 N18726 0 diode
R18727 N18726 N18727 10
D18727 N18727 0 diode
R18728 N18727 N18728 10
D18728 N18728 0 diode
R18729 N18728 N18729 10
D18729 N18729 0 diode
R18730 N18729 N18730 10
D18730 N18730 0 diode
R18731 N18730 N18731 10
D18731 N18731 0 diode
R18732 N18731 N18732 10
D18732 N18732 0 diode
R18733 N18732 N18733 10
D18733 N18733 0 diode
R18734 N18733 N18734 10
D18734 N18734 0 diode
R18735 N18734 N18735 10
D18735 N18735 0 diode
R18736 N18735 N18736 10
D18736 N18736 0 diode
R18737 N18736 N18737 10
D18737 N18737 0 diode
R18738 N18737 N18738 10
D18738 N18738 0 diode
R18739 N18738 N18739 10
D18739 N18739 0 diode
R18740 N18739 N18740 10
D18740 N18740 0 diode
R18741 N18740 N18741 10
D18741 N18741 0 diode
R18742 N18741 N18742 10
D18742 N18742 0 diode
R18743 N18742 N18743 10
D18743 N18743 0 diode
R18744 N18743 N18744 10
D18744 N18744 0 diode
R18745 N18744 N18745 10
D18745 N18745 0 diode
R18746 N18745 N18746 10
D18746 N18746 0 diode
R18747 N18746 N18747 10
D18747 N18747 0 diode
R18748 N18747 N18748 10
D18748 N18748 0 diode
R18749 N18748 N18749 10
D18749 N18749 0 diode
R18750 N18749 N18750 10
D18750 N18750 0 diode
R18751 N18750 N18751 10
D18751 N18751 0 diode
R18752 N18751 N18752 10
D18752 N18752 0 diode
R18753 N18752 N18753 10
D18753 N18753 0 diode
R18754 N18753 N18754 10
D18754 N18754 0 diode
R18755 N18754 N18755 10
D18755 N18755 0 diode
R18756 N18755 N18756 10
D18756 N18756 0 diode
R18757 N18756 N18757 10
D18757 N18757 0 diode
R18758 N18757 N18758 10
D18758 N18758 0 diode
R18759 N18758 N18759 10
D18759 N18759 0 diode
R18760 N18759 N18760 10
D18760 N18760 0 diode
R18761 N18760 N18761 10
D18761 N18761 0 diode
R18762 N18761 N18762 10
D18762 N18762 0 diode
R18763 N18762 N18763 10
D18763 N18763 0 diode
R18764 N18763 N18764 10
D18764 N18764 0 diode
R18765 N18764 N18765 10
D18765 N18765 0 diode
R18766 N18765 N18766 10
D18766 N18766 0 diode
R18767 N18766 N18767 10
D18767 N18767 0 diode
R18768 N18767 N18768 10
D18768 N18768 0 diode
R18769 N18768 N18769 10
D18769 N18769 0 diode
R18770 N18769 N18770 10
D18770 N18770 0 diode
R18771 N18770 N18771 10
D18771 N18771 0 diode
R18772 N18771 N18772 10
D18772 N18772 0 diode
R18773 N18772 N18773 10
D18773 N18773 0 diode
R18774 N18773 N18774 10
D18774 N18774 0 diode
R18775 N18774 N18775 10
D18775 N18775 0 diode
R18776 N18775 N18776 10
D18776 N18776 0 diode
R18777 N18776 N18777 10
D18777 N18777 0 diode
R18778 N18777 N18778 10
D18778 N18778 0 diode
R18779 N18778 N18779 10
D18779 N18779 0 diode
R18780 N18779 N18780 10
D18780 N18780 0 diode
R18781 N18780 N18781 10
D18781 N18781 0 diode
R18782 N18781 N18782 10
D18782 N18782 0 diode
R18783 N18782 N18783 10
D18783 N18783 0 diode
R18784 N18783 N18784 10
D18784 N18784 0 diode
R18785 N18784 N18785 10
D18785 N18785 0 diode
R18786 N18785 N18786 10
D18786 N18786 0 diode
R18787 N18786 N18787 10
D18787 N18787 0 diode
R18788 N18787 N18788 10
D18788 N18788 0 diode
R18789 N18788 N18789 10
D18789 N18789 0 diode
R18790 N18789 N18790 10
D18790 N18790 0 diode
R18791 N18790 N18791 10
D18791 N18791 0 diode
R18792 N18791 N18792 10
D18792 N18792 0 diode
R18793 N18792 N18793 10
D18793 N18793 0 diode
R18794 N18793 N18794 10
D18794 N18794 0 diode
R18795 N18794 N18795 10
D18795 N18795 0 diode
R18796 N18795 N18796 10
D18796 N18796 0 diode
R18797 N18796 N18797 10
D18797 N18797 0 diode
R18798 N18797 N18798 10
D18798 N18798 0 diode
R18799 N18798 N18799 10
D18799 N18799 0 diode
R18800 N18799 N18800 10
D18800 N18800 0 diode
R18801 N18800 N18801 10
D18801 N18801 0 diode
R18802 N18801 N18802 10
D18802 N18802 0 diode
R18803 N18802 N18803 10
D18803 N18803 0 diode
R18804 N18803 N18804 10
D18804 N18804 0 diode
R18805 N18804 N18805 10
D18805 N18805 0 diode
R18806 N18805 N18806 10
D18806 N18806 0 diode
R18807 N18806 N18807 10
D18807 N18807 0 diode
R18808 N18807 N18808 10
D18808 N18808 0 diode
R18809 N18808 N18809 10
D18809 N18809 0 diode
R18810 N18809 N18810 10
D18810 N18810 0 diode
R18811 N18810 N18811 10
D18811 N18811 0 diode
R18812 N18811 N18812 10
D18812 N18812 0 diode
R18813 N18812 N18813 10
D18813 N18813 0 diode
R18814 N18813 N18814 10
D18814 N18814 0 diode
R18815 N18814 N18815 10
D18815 N18815 0 diode
R18816 N18815 N18816 10
D18816 N18816 0 diode
R18817 N18816 N18817 10
D18817 N18817 0 diode
R18818 N18817 N18818 10
D18818 N18818 0 diode
R18819 N18818 N18819 10
D18819 N18819 0 diode
R18820 N18819 N18820 10
D18820 N18820 0 diode
R18821 N18820 N18821 10
D18821 N18821 0 diode
R18822 N18821 N18822 10
D18822 N18822 0 diode
R18823 N18822 N18823 10
D18823 N18823 0 diode
R18824 N18823 N18824 10
D18824 N18824 0 diode
R18825 N18824 N18825 10
D18825 N18825 0 diode
R18826 N18825 N18826 10
D18826 N18826 0 diode
R18827 N18826 N18827 10
D18827 N18827 0 diode
R18828 N18827 N18828 10
D18828 N18828 0 diode
R18829 N18828 N18829 10
D18829 N18829 0 diode
R18830 N18829 N18830 10
D18830 N18830 0 diode
R18831 N18830 N18831 10
D18831 N18831 0 diode
R18832 N18831 N18832 10
D18832 N18832 0 diode
R18833 N18832 N18833 10
D18833 N18833 0 diode
R18834 N18833 N18834 10
D18834 N18834 0 diode
R18835 N18834 N18835 10
D18835 N18835 0 diode
R18836 N18835 N18836 10
D18836 N18836 0 diode
R18837 N18836 N18837 10
D18837 N18837 0 diode
R18838 N18837 N18838 10
D18838 N18838 0 diode
R18839 N18838 N18839 10
D18839 N18839 0 diode
R18840 N18839 N18840 10
D18840 N18840 0 diode
R18841 N18840 N18841 10
D18841 N18841 0 diode
R18842 N18841 N18842 10
D18842 N18842 0 diode
R18843 N18842 N18843 10
D18843 N18843 0 diode
R18844 N18843 N18844 10
D18844 N18844 0 diode
R18845 N18844 N18845 10
D18845 N18845 0 diode
R18846 N18845 N18846 10
D18846 N18846 0 diode
R18847 N18846 N18847 10
D18847 N18847 0 diode
R18848 N18847 N18848 10
D18848 N18848 0 diode
R18849 N18848 N18849 10
D18849 N18849 0 diode
R18850 N18849 N18850 10
D18850 N18850 0 diode
R18851 N18850 N18851 10
D18851 N18851 0 diode
R18852 N18851 N18852 10
D18852 N18852 0 diode
R18853 N18852 N18853 10
D18853 N18853 0 diode
R18854 N18853 N18854 10
D18854 N18854 0 diode
R18855 N18854 N18855 10
D18855 N18855 0 diode
R18856 N18855 N18856 10
D18856 N18856 0 diode
R18857 N18856 N18857 10
D18857 N18857 0 diode
R18858 N18857 N18858 10
D18858 N18858 0 diode
R18859 N18858 N18859 10
D18859 N18859 0 diode
R18860 N18859 N18860 10
D18860 N18860 0 diode
R18861 N18860 N18861 10
D18861 N18861 0 diode
R18862 N18861 N18862 10
D18862 N18862 0 diode
R18863 N18862 N18863 10
D18863 N18863 0 diode
R18864 N18863 N18864 10
D18864 N18864 0 diode
R18865 N18864 N18865 10
D18865 N18865 0 diode
R18866 N18865 N18866 10
D18866 N18866 0 diode
R18867 N18866 N18867 10
D18867 N18867 0 diode
R18868 N18867 N18868 10
D18868 N18868 0 diode
R18869 N18868 N18869 10
D18869 N18869 0 diode
R18870 N18869 N18870 10
D18870 N18870 0 diode
R18871 N18870 N18871 10
D18871 N18871 0 diode
R18872 N18871 N18872 10
D18872 N18872 0 diode
R18873 N18872 N18873 10
D18873 N18873 0 diode
R18874 N18873 N18874 10
D18874 N18874 0 diode
R18875 N18874 N18875 10
D18875 N18875 0 diode
R18876 N18875 N18876 10
D18876 N18876 0 diode
R18877 N18876 N18877 10
D18877 N18877 0 diode
R18878 N18877 N18878 10
D18878 N18878 0 diode
R18879 N18878 N18879 10
D18879 N18879 0 diode
R18880 N18879 N18880 10
D18880 N18880 0 diode
R18881 N18880 N18881 10
D18881 N18881 0 diode
R18882 N18881 N18882 10
D18882 N18882 0 diode
R18883 N18882 N18883 10
D18883 N18883 0 diode
R18884 N18883 N18884 10
D18884 N18884 0 diode
R18885 N18884 N18885 10
D18885 N18885 0 diode
R18886 N18885 N18886 10
D18886 N18886 0 diode
R18887 N18886 N18887 10
D18887 N18887 0 diode
R18888 N18887 N18888 10
D18888 N18888 0 diode
R18889 N18888 N18889 10
D18889 N18889 0 diode
R18890 N18889 N18890 10
D18890 N18890 0 diode
R18891 N18890 N18891 10
D18891 N18891 0 diode
R18892 N18891 N18892 10
D18892 N18892 0 diode
R18893 N18892 N18893 10
D18893 N18893 0 diode
R18894 N18893 N18894 10
D18894 N18894 0 diode
R18895 N18894 N18895 10
D18895 N18895 0 diode
R18896 N18895 N18896 10
D18896 N18896 0 diode
R18897 N18896 N18897 10
D18897 N18897 0 diode
R18898 N18897 N18898 10
D18898 N18898 0 diode
R18899 N18898 N18899 10
D18899 N18899 0 diode
R18900 N18899 N18900 10
D18900 N18900 0 diode
R18901 N18900 N18901 10
D18901 N18901 0 diode
R18902 N18901 N18902 10
D18902 N18902 0 diode
R18903 N18902 N18903 10
D18903 N18903 0 diode
R18904 N18903 N18904 10
D18904 N18904 0 diode
R18905 N18904 N18905 10
D18905 N18905 0 diode
R18906 N18905 N18906 10
D18906 N18906 0 diode
R18907 N18906 N18907 10
D18907 N18907 0 diode
R18908 N18907 N18908 10
D18908 N18908 0 diode
R18909 N18908 N18909 10
D18909 N18909 0 diode
R18910 N18909 N18910 10
D18910 N18910 0 diode
R18911 N18910 N18911 10
D18911 N18911 0 diode
R18912 N18911 N18912 10
D18912 N18912 0 diode
R18913 N18912 N18913 10
D18913 N18913 0 diode
R18914 N18913 N18914 10
D18914 N18914 0 diode
R18915 N18914 N18915 10
D18915 N18915 0 diode
R18916 N18915 N18916 10
D18916 N18916 0 diode
R18917 N18916 N18917 10
D18917 N18917 0 diode
R18918 N18917 N18918 10
D18918 N18918 0 diode
R18919 N18918 N18919 10
D18919 N18919 0 diode
R18920 N18919 N18920 10
D18920 N18920 0 diode
R18921 N18920 N18921 10
D18921 N18921 0 diode
R18922 N18921 N18922 10
D18922 N18922 0 diode
R18923 N18922 N18923 10
D18923 N18923 0 diode
R18924 N18923 N18924 10
D18924 N18924 0 diode
R18925 N18924 N18925 10
D18925 N18925 0 diode
R18926 N18925 N18926 10
D18926 N18926 0 diode
R18927 N18926 N18927 10
D18927 N18927 0 diode
R18928 N18927 N18928 10
D18928 N18928 0 diode
R18929 N18928 N18929 10
D18929 N18929 0 diode
R18930 N18929 N18930 10
D18930 N18930 0 diode
R18931 N18930 N18931 10
D18931 N18931 0 diode
R18932 N18931 N18932 10
D18932 N18932 0 diode
R18933 N18932 N18933 10
D18933 N18933 0 diode
R18934 N18933 N18934 10
D18934 N18934 0 diode
R18935 N18934 N18935 10
D18935 N18935 0 diode
R18936 N18935 N18936 10
D18936 N18936 0 diode
R18937 N18936 N18937 10
D18937 N18937 0 diode
R18938 N18937 N18938 10
D18938 N18938 0 diode
R18939 N18938 N18939 10
D18939 N18939 0 diode
R18940 N18939 N18940 10
D18940 N18940 0 diode
R18941 N18940 N18941 10
D18941 N18941 0 diode
R18942 N18941 N18942 10
D18942 N18942 0 diode
R18943 N18942 N18943 10
D18943 N18943 0 diode
R18944 N18943 N18944 10
D18944 N18944 0 diode
R18945 N18944 N18945 10
D18945 N18945 0 diode
R18946 N18945 N18946 10
D18946 N18946 0 diode
R18947 N18946 N18947 10
D18947 N18947 0 diode
R18948 N18947 N18948 10
D18948 N18948 0 diode
R18949 N18948 N18949 10
D18949 N18949 0 diode
R18950 N18949 N18950 10
D18950 N18950 0 diode
R18951 N18950 N18951 10
D18951 N18951 0 diode
R18952 N18951 N18952 10
D18952 N18952 0 diode
R18953 N18952 N18953 10
D18953 N18953 0 diode
R18954 N18953 N18954 10
D18954 N18954 0 diode
R18955 N18954 N18955 10
D18955 N18955 0 diode
R18956 N18955 N18956 10
D18956 N18956 0 diode
R18957 N18956 N18957 10
D18957 N18957 0 diode
R18958 N18957 N18958 10
D18958 N18958 0 diode
R18959 N18958 N18959 10
D18959 N18959 0 diode
R18960 N18959 N18960 10
D18960 N18960 0 diode
R18961 N18960 N18961 10
D18961 N18961 0 diode
R18962 N18961 N18962 10
D18962 N18962 0 diode
R18963 N18962 N18963 10
D18963 N18963 0 diode
R18964 N18963 N18964 10
D18964 N18964 0 diode
R18965 N18964 N18965 10
D18965 N18965 0 diode
R18966 N18965 N18966 10
D18966 N18966 0 diode
R18967 N18966 N18967 10
D18967 N18967 0 diode
R18968 N18967 N18968 10
D18968 N18968 0 diode
R18969 N18968 N18969 10
D18969 N18969 0 diode
R18970 N18969 N18970 10
D18970 N18970 0 diode
R18971 N18970 N18971 10
D18971 N18971 0 diode
R18972 N18971 N18972 10
D18972 N18972 0 diode
R18973 N18972 N18973 10
D18973 N18973 0 diode
R18974 N18973 N18974 10
D18974 N18974 0 diode
R18975 N18974 N18975 10
D18975 N18975 0 diode
R18976 N18975 N18976 10
D18976 N18976 0 diode
R18977 N18976 N18977 10
D18977 N18977 0 diode
R18978 N18977 N18978 10
D18978 N18978 0 diode
R18979 N18978 N18979 10
D18979 N18979 0 diode
R18980 N18979 N18980 10
D18980 N18980 0 diode
R18981 N18980 N18981 10
D18981 N18981 0 diode
R18982 N18981 N18982 10
D18982 N18982 0 diode
R18983 N18982 N18983 10
D18983 N18983 0 diode
R18984 N18983 N18984 10
D18984 N18984 0 diode
R18985 N18984 N18985 10
D18985 N18985 0 diode
R18986 N18985 N18986 10
D18986 N18986 0 diode
R18987 N18986 N18987 10
D18987 N18987 0 diode
R18988 N18987 N18988 10
D18988 N18988 0 diode
R18989 N18988 N18989 10
D18989 N18989 0 diode
R18990 N18989 N18990 10
D18990 N18990 0 diode
R18991 N18990 N18991 10
D18991 N18991 0 diode
R18992 N18991 N18992 10
D18992 N18992 0 diode
R18993 N18992 N18993 10
D18993 N18993 0 diode
R18994 N18993 N18994 10
D18994 N18994 0 diode
R18995 N18994 N18995 10
D18995 N18995 0 diode
R18996 N18995 N18996 10
D18996 N18996 0 diode
R18997 N18996 N18997 10
D18997 N18997 0 diode
R18998 N18997 N18998 10
D18998 N18998 0 diode
R18999 N18998 N18999 10
D18999 N18999 0 diode
R19000 N18999 N19000 10
D19000 N19000 0 diode
R19001 N19000 N19001 10
D19001 N19001 0 diode
R19002 N19001 N19002 10
D19002 N19002 0 diode
R19003 N19002 N19003 10
D19003 N19003 0 diode
R19004 N19003 N19004 10
D19004 N19004 0 diode
R19005 N19004 N19005 10
D19005 N19005 0 diode
R19006 N19005 N19006 10
D19006 N19006 0 diode
R19007 N19006 N19007 10
D19007 N19007 0 diode
R19008 N19007 N19008 10
D19008 N19008 0 diode
R19009 N19008 N19009 10
D19009 N19009 0 diode
R19010 N19009 N19010 10
D19010 N19010 0 diode
R19011 N19010 N19011 10
D19011 N19011 0 diode
R19012 N19011 N19012 10
D19012 N19012 0 diode
R19013 N19012 N19013 10
D19013 N19013 0 diode
R19014 N19013 N19014 10
D19014 N19014 0 diode
R19015 N19014 N19015 10
D19015 N19015 0 diode
R19016 N19015 N19016 10
D19016 N19016 0 diode
R19017 N19016 N19017 10
D19017 N19017 0 diode
R19018 N19017 N19018 10
D19018 N19018 0 diode
R19019 N19018 N19019 10
D19019 N19019 0 diode
R19020 N19019 N19020 10
D19020 N19020 0 diode
R19021 N19020 N19021 10
D19021 N19021 0 diode
R19022 N19021 N19022 10
D19022 N19022 0 diode
R19023 N19022 N19023 10
D19023 N19023 0 diode
R19024 N19023 N19024 10
D19024 N19024 0 diode
R19025 N19024 N19025 10
D19025 N19025 0 diode
R19026 N19025 N19026 10
D19026 N19026 0 diode
R19027 N19026 N19027 10
D19027 N19027 0 diode
R19028 N19027 N19028 10
D19028 N19028 0 diode
R19029 N19028 N19029 10
D19029 N19029 0 diode
R19030 N19029 N19030 10
D19030 N19030 0 diode
R19031 N19030 N19031 10
D19031 N19031 0 diode
R19032 N19031 N19032 10
D19032 N19032 0 diode
R19033 N19032 N19033 10
D19033 N19033 0 diode
R19034 N19033 N19034 10
D19034 N19034 0 diode
R19035 N19034 N19035 10
D19035 N19035 0 diode
R19036 N19035 N19036 10
D19036 N19036 0 diode
R19037 N19036 N19037 10
D19037 N19037 0 diode
R19038 N19037 N19038 10
D19038 N19038 0 diode
R19039 N19038 N19039 10
D19039 N19039 0 diode
R19040 N19039 N19040 10
D19040 N19040 0 diode
R19041 N19040 N19041 10
D19041 N19041 0 diode
R19042 N19041 N19042 10
D19042 N19042 0 diode
R19043 N19042 N19043 10
D19043 N19043 0 diode
R19044 N19043 N19044 10
D19044 N19044 0 diode
R19045 N19044 N19045 10
D19045 N19045 0 diode
R19046 N19045 N19046 10
D19046 N19046 0 diode
R19047 N19046 N19047 10
D19047 N19047 0 diode
R19048 N19047 N19048 10
D19048 N19048 0 diode
R19049 N19048 N19049 10
D19049 N19049 0 diode
R19050 N19049 N19050 10
D19050 N19050 0 diode
R19051 N19050 N19051 10
D19051 N19051 0 diode
R19052 N19051 N19052 10
D19052 N19052 0 diode
R19053 N19052 N19053 10
D19053 N19053 0 diode
R19054 N19053 N19054 10
D19054 N19054 0 diode
R19055 N19054 N19055 10
D19055 N19055 0 diode
R19056 N19055 N19056 10
D19056 N19056 0 diode
R19057 N19056 N19057 10
D19057 N19057 0 diode
R19058 N19057 N19058 10
D19058 N19058 0 diode
R19059 N19058 N19059 10
D19059 N19059 0 diode
R19060 N19059 N19060 10
D19060 N19060 0 diode
R19061 N19060 N19061 10
D19061 N19061 0 diode
R19062 N19061 N19062 10
D19062 N19062 0 diode
R19063 N19062 N19063 10
D19063 N19063 0 diode
R19064 N19063 N19064 10
D19064 N19064 0 diode
R19065 N19064 N19065 10
D19065 N19065 0 diode
R19066 N19065 N19066 10
D19066 N19066 0 diode
R19067 N19066 N19067 10
D19067 N19067 0 diode
R19068 N19067 N19068 10
D19068 N19068 0 diode
R19069 N19068 N19069 10
D19069 N19069 0 diode
R19070 N19069 N19070 10
D19070 N19070 0 diode
R19071 N19070 N19071 10
D19071 N19071 0 diode
R19072 N19071 N19072 10
D19072 N19072 0 diode
R19073 N19072 N19073 10
D19073 N19073 0 diode
R19074 N19073 N19074 10
D19074 N19074 0 diode
R19075 N19074 N19075 10
D19075 N19075 0 diode
R19076 N19075 N19076 10
D19076 N19076 0 diode
R19077 N19076 N19077 10
D19077 N19077 0 diode
R19078 N19077 N19078 10
D19078 N19078 0 diode
R19079 N19078 N19079 10
D19079 N19079 0 diode
R19080 N19079 N19080 10
D19080 N19080 0 diode
R19081 N19080 N19081 10
D19081 N19081 0 diode
R19082 N19081 N19082 10
D19082 N19082 0 diode
R19083 N19082 N19083 10
D19083 N19083 0 diode
R19084 N19083 N19084 10
D19084 N19084 0 diode
R19085 N19084 N19085 10
D19085 N19085 0 diode
R19086 N19085 N19086 10
D19086 N19086 0 diode
R19087 N19086 N19087 10
D19087 N19087 0 diode
R19088 N19087 N19088 10
D19088 N19088 0 diode
R19089 N19088 N19089 10
D19089 N19089 0 diode
R19090 N19089 N19090 10
D19090 N19090 0 diode
R19091 N19090 N19091 10
D19091 N19091 0 diode
R19092 N19091 N19092 10
D19092 N19092 0 diode
R19093 N19092 N19093 10
D19093 N19093 0 diode
R19094 N19093 N19094 10
D19094 N19094 0 diode
R19095 N19094 N19095 10
D19095 N19095 0 diode
R19096 N19095 N19096 10
D19096 N19096 0 diode
R19097 N19096 N19097 10
D19097 N19097 0 diode
R19098 N19097 N19098 10
D19098 N19098 0 diode
R19099 N19098 N19099 10
D19099 N19099 0 diode
R19100 N19099 N19100 10
D19100 N19100 0 diode
R19101 N19100 N19101 10
D19101 N19101 0 diode
R19102 N19101 N19102 10
D19102 N19102 0 diode
R19103 N19102 N19103 10
D19103 N19103 0 diode
R19104 N19103 N19104 10
D19104 N19104 0 diode
R19105 N19104 N19105 10
D19105 N19105 0 diode
R19106 N19105 N19106 10
D19106 N19106 0 diode
R19107 N19106 N19107 10
D19107 N19107 0 diode
R19108 N19107 N19108 10
D19108 N19108 0 diode
R19109 N19108 N19109 10
D19109 N19109 0 diode
R19110 N19109 N19110 10
D19110 N19110 0 diode
R19111 N19110 N19111 10
D19111 N19111 0 diode
R19112 N19111 N19112 10
D19112 N19112 0 diode
R19113 N19112 N19113 10
D19113 N19113 0 diode
R19114 N19113 N19114 10
D19114 N19114 0 diode
R19115 N19114 N19115 10
D19115 N19115 0 diode
R19116 N19115 N19116 10
D19116 N19116 0 diode
R19117 N19116 N19117 10
D19117 N19117 0 diode
R19118 N19117 N19118 10
D19118 N19118 0 diode
R19119 N19118 N19119 10
D19119 N19119 0 diode
R19120 N19119 N19120 10
D19120 N19120 0 diode
R19121 N19120 N19121 10
D19121 N19121 0 diode
R19122 N19121 N19122 10
D19122 N19122 0 diode
R19123 N19122 N19123 10
D19123 N19123 0 diode
R19124 N19123 N19124 10
D19124 N19124 0 diode
R19125 N19124 N19125 10
D19125 N19125 0 diode
R19126 N19125 N19126 10
D19126 N19126 0 diode
R19127 N19126 N19127 10
D19127 N19127 0 diode
R19128 N19127 N19128 10
D19128 N19128 0 diode
R19129 N19128 N19129 10
D19129 N19129 0 diode
R19130 N19129 N19130 10
D19130 N19130 0 diode
R19131 N19130 N19131 10
D19131 N19131 0 diode
R19132 N19131 N19132 10
D19132 N19132 0 diode
R19133 N19132 N19133 10
D19133 N19133 0 diode
R19134 N19133 N19134 10
D19134 N19134 0 diode
R19135 N19134 N19135 10
D19135 N19135 0 diode
R19136 N19135 N19136 10
D19136 N19136 0 diode
R19137 N19136 N19137 10
D19137 N19137 0 diode
R19138 N19137 N19138 10
D19138 N19138 0 diode
R19139 N19138 N19139 10
D19139 N19139 0 diode
R19140 N19139 N19140 10
D19140 N19140 0 diode
R19141 N19140 N19141 10
D19141 N19141 0 diode
R19142 N19141 N19142 10
D19142 N19142 0 diode
R19143 N19142 N19143 10
D19143 N19143 0 diode
R19144 N19143 N19144 10
D19144 N19144 0 diode
R19145 N19144 N19145 10
D19145 N19145 0 diode
R19146 N19145 N19146 10
D19146 N19146 0 diode
R19147 N19146 N19147 10
D19147 N19147 0 diode
R19148 N19147 N19148 10
D19148 N19148 0 diode
R19149 N19148 N19149 10
D19149 N19149 0 diode
R19150 N19149 N19150 10
D19150 N19150 0 diode
R19151 N19150 N19151 10
D19151 N19151 0 diode
R19152 N19151 N19152 10
D19152 N19152 0 diode
R19153 N19152 N19153 10
D19153 N19153 0 diode
R19154 N19153 N19154 10
D19154 N19154 0 diode
R19155 N19154 N19155 10
D19155 N19155 0 diode
R19156 N19155 N19156 10
D19156 N19156 0 diode
R19157 N19156 N19157 10
D19157 N19157 0 diode
R19158 N19157 N19158 10
D19158 N19158 0 diode
R19159 N19158 N19159 10
D19159 N19159 0 diode
R19160 N19159 N19160 10
D19160 N19160 0 diode
R19161 N19160 N19161 10
D19161 N19161 0 diode
R19162 N19161 N19162 10
D19162 N19162 0 diode
R19163 N19162 N19163 10
D19163 N19163 0 diode
R19164 N19163 N19164 10
D19164 N19164 0 diode
R19165 N19164 N19165 10
D19165 N19165 0 diode
R19166 N19165 N19166 10
D19166 N19166 0 diode
R19167 N19166 N19167 10
D19167 N19167 0 diode
R19168 N19167 N19168 10
D19168 N19168 0 diode
R19169 N19168 N19169 10
D19169 N19169 0 diode
R19170 N19169 N19170 10
D19170 N19170 0 diode
R19171 N19170 N19171 10
D19171 N19171 0 diode
R19172 N19171 N19172 10
D19172 N19172 0 diode
R19173 N19172 N19173 10
D19173 N19173 0 diode
R19174 N19173 N19174 10
D19174 N19174 0 diode
R19175 N19174 N19175 10
D19175 N19175 0 diode
R19176 N19175 N19176 10
D19176 N19176 0 diode
R19177 N19176 N19177 10
D19177 N19177 0 diode
R19178 N19177 N19178 10
D19178 N19178 0 diode
R19179 N19178 N19179 10
D19179 N19179 0 diode
R19180 N19179 N19180 10
D19180 N19180 0 diode
R19181 N19180 N19181 10
D19181 N19181 0 diode
R19182 N19181 N19182 10
D19182 N19182 0 diode
R19183 N19182 N19183 10
D19183 N19183 0 diode
R19184 N19183 N19184 10
D19184 N19184 0 diode
R19185 N19184 N19185 10
D19185 N19185 0 diode
R19186 N19185 N19186 10
D19186 N19186 0 diode
R19187 N19186 N19187 10
D19187 N19187 0 diode
R19188 N19187 N19188 10
D19188 N19188 0 diode
R19189 N19188 N19189 10
D19189 N19189 0 diode
R19190 N19189 N19190 10
D19190 N19190 0 diode
R19191 N19190 N19191 10
D19191 N19191 0 diode
R19192 N19191 N19192 10
D19192 N19192 0 diode
R19193 N19192 N19193 10
D19193 N19193 0 diode
R19194 N19193 N19194 10
D19194 N19194 0 diode
R19195 N19194 N19195 10
D19195 N19195 0 diode
R19196 N19195 N19196 10
D19196 N19196 0 diode
R19197 N19196 N19197 10
D19197 N19197 0 diode
R19198 N19197 N19198 10
D19198 N19198 0 diode
R19199 N19198 N19199 10
D19199 N19199 0 diode
R19200 N19199 N19200 10
D19200 N19200 0 diode
R19201 N19200 N19201 10
D19201 N19201 0 diode
R19202 N19201 N19202 10
D19202 N19202 0 diode
R19203 N19202 N19203 10
D19203 N19203 0 diode
R19204 N19203 N19204 10
D19204 N19204 0 diode
R19205 N19204 N19205 10
D19205 N19205 0 diode
R19206 N19205 N19206 10
D19206 N19206 0 diode
R19207 N19206 N19207 10
D19207 N19207 0 diode
R19208 N19207 N19208 10
D19208 N19208 0 diode
R19209 N19208 N19209 10
D19209 N19209 0 diode
R19210 N19209 N19210 10
D19210 N19210 0 diode
R19211 N19210 N19211 10
D19211 N19211 0 diode
R19212 N19211 N19212 10
D19212 N19212 0 diode
R19213 N19212 N19213 10
D19213 N19213 0 diode
R19214 N19213 N19214 10
D19214 N19214 0 diode
R19215 N19214 N19215 10
D19215 N19215 0 diode
R19216 N19215 N19216 10
D19216 N19216 0 diode
R19217 N19216 N19217 10
D19217 N19217 0 diode
R19218 N19217 N19218 10
D19218 N19218 0 diode
R19219 N19218 N19219 10
D19219 N19219 0 diode
R19220 N19219 N19220 10
D19220 N19220 0 diode
R19221 N19220 N19221 10
D19221 N19221 0 diode
R19222 N19221 N19222 10
D19222 N19222 0 diode
R19223 N19222 N19223 10
D19223 N19223 0 diode
R19224 N19223 N19224 10
D19224 N19224 0 diode
R19225 N19224 N19225 10
D19225 N19225 0 diode
R19226 N19225 N19226 10
D19226 N19226 0 diode
R19227 N19226 N19227 10
D19227 N19227 0 diode
R19228 N19227 N19228 10
D19228 N19228 0 diode
R19229 N19228 N19229 10
D19229 N19229 0 diode
R19230 N19229 N19230 10
D19230 N19230 0 diode
R19231 N19230 N19231 10
D19231 N19231 0 diode
R19232 N19231 N19232 10
D19232 N19232 0 diode
R19233 N19232 N19233 10
D19233 N19233 0 diode
R19234 N19233 N19234 10
D19234 N19234 0 diode
R19235 N19234 N19235 10
D19235 N19235 0 diode
R19236 N19235 N19236 10
D19236 N19236 0 diode
R19237 N19236 N19237 10
D19237 N19237 0 diode
R19238 N19237 N19238 10
D19238 N19238 0 diode
R19239 N19238 N19239 10
D19239 N19239 0 diode
R19240 N19239 N19240 10
D19240 N19240 0 diode
R19241 N19240 N19241 10
D19241 N19241 0 diode
R19242 N19241 N19242 10
D19242 N19242 0 diode
R19243 N19242 N19243 10
D19243 N19243 0 diode
R19244 N19243 N19244 10
D19244 N19244 0 diode
R19245 N19244 N19245 10
D19245 N19245 0 diode
R19246 N19245 N19246 10
D19246 N19246 0 diode
R19247 N19246 N19247 10
D19247 N19247 0 diode
R19248 N19247 N19248 10
D19248 N19248 0 diode
R19249 N19248 N19249 10
D19249 N19249 0 diode
R19250 N19249 N19250 10
D19250 N19250 0 diode
R19251 N19250 N19251 10
D19251 N19251 0 diode
R19252 N19251 N19252 10
D19252 N19252 0 diode
R19253 N19252 N19253 10
D19253 N19253 0 diode
R19254 N19253 N19254 10
D19254 N19254 0 diode
R19255 N19254 N19255 10
D19255 N19255 0 diode
R19256 N19255 N19256 10
D19256 N19256 0 diode
R19257 N19256 N19257 10
D19257 N19257 0 diode
R19258 N19257 N19258 10
D19258 N19258 0 diode
R19259 N19258 N19259 10
D19259 N19259 0 diode
R19260 N19259 N19260 10
D19260 N19260 0 diode
R19261 N19260 N19261 10
D19261 N19261 0 diode
R19262 N19261 N19262 10
D19262 N19262 0 diode
R19263 N19262 N19263 10
D19263 N19263 0 diode
R19264 N19263 N19264 10
D19264 N19264 0 diode
R19265 N19264 N19265 10
D19265 N19265 0 diode
R19266 N19265 N19266 10
D19266 N19266 0 diode
R19267 N19266 N19267 10
D19267 N19267 0 diode
R19268 N19267 N19268 10
D19268 N19268 0 diode
R19269 N19268 N19269 10
D19269 N19269 0 diode
R19270 N19269 N19270 10
D19270 N19270 0 diode
R19271 N19270 N19271 10
D19271 N19271 0 diode
R19272 N19271 N19272 10
D19272 N19272 0 diode
R19273 N19272 N19273 10
D19273 N19273 0 diode
R19274 N19273 N19274 10
D19274 N19274 0 diode
R19275 N19274 N19275 10
D19275 N19275 0 diode
R19276 N19275 N19276 10
D19276 N19276 0 diode
R19277 N19276 N19277 10
D19277 N19277 0 diode
R19278 N19277 N19278 10
D19278 N19278 0 diode
R19279 N19278 N19279 10
D19279 N19279 0 diode
R19280 N19279 N19280 10
D19280 N19280 0 diode
R19281 N19280 N19281 10
D19281 N19281 0 diode
R19282 N19281 N19282 10
D19282 N19282 0 diode
R19283 N19282 N19283 10
D19283 N19283 0 diode
R19284 N19283 N19284 10
D19284 N19284 0 diode
R19285 N19284 N19285 10
D19285 N19285 0 diode
R19286 N19285 N19286 10
D19286 N19286 0 diode
R19287 N19286 N19287 10
D19287 N19287 0 diode
R19288 N19287 N19288 10
D19288 N19288 0 diode
R19289 N19288 N19289 10
D19289 N19289 0 diode
R19290 N19289 N19290 10
D19290 N19290 0 diode
R19291 N19290 N19291 10
D19291 N19291 0 diode
R19292 N19291 N19292 10
D19292 N19292 0 diode
R19293 N19292 N19293 10
D19293 N19293 0 diode
R19294 N19293 N19294 10
D19294 N19294 0 diode
R19295 N19294 N19295 10
D19295 N19295 0 diode
R19296 N19295 N19296 10
D19296 N19296 0 diode
R19297 N19296 N19297 10
D19297 N19297 0 diode
R19298 N19297 N19298 10
D19298 N19298 0 diode
R19299 N19298 N19299 10
D19299 N19299 0 diode
R19300 N19299 N19300 10
D19300 N19300 0 diode
R19301 N19300 N19301 10
D19301 N19301 0 diode
R19302 N19301 N19302 10
D19302 N19302 0 diode
R19303 N19302 N19303 10
D19303 N19303 0 diode
R19304 N19303 N19304 10
D19304 N19304 0 diode
R19305 N19304 N19305 10
D19305 N19305 0 diode
R19306 N19305 N19306 10
D19306 N19306 0 diode
R19307 N19306 N19307 10
D19307 N19307 0 diode
R19308 N19307 N19308 10
D19308 N19308 0 diode
R19309 N19308 N19309 10
D19309 N19309 0 diode
R19310 N19309 N19310 10
D19310 N19310 0 diode
R19311 N19310 N19311 10
D19311 N19311 0 diode
R19312 N19311 N19312 10
D19312 N19312 0 diode
R19313 N19312 N19313 10
D19313 N19313 0 diode
R19314 N19313 N19314 10
D19314 N19314 0 diode
R19315 N19314 N19315 10
D19315 N19315 0 diode
R19316 N19315 N19316 10
D19316 N19316 0 diode
R19317 N19316 N19317 10
D19317 N19317 0 diode
R19318 N19317 N19318 10
D19318 N19318 0 diode
R19319 N19318 N19319 10
D19319 N19319 0 diode
R19320 N19319 N19320 10
D19320 N19320 0 diode
R19321 N19320 N19321 10
D19321 N19321 0 diode
R19322 N19321 N19322 10
D19322 N19322 0 diode
R19323 N19322 N19323 10
D19323 N19323 0 diode
R19324 N19323 N19324 10
D19324 N19324 0 diode
R19325 N19324 N19325 10
D19325 N19325 0 diode
R19326 N19325 N19326 10
D19326 N19326 0 diode
R19327 N19326 N19327 10
D19327 N19327 0 diode
R19328 N19327 N19328 10
D19328 N19328 0 diode
R19329 N19328 N19329 10
D19329 N19329 0 diode
R19330 N19329 N19330 10
D19330 N19330 0 diode
R19331 N19330 N19331 10
D19331 N19331 0 diode
R19332 N19331 N19332 10
D19332 N19332 0 diode
R19333 N19332 N19333 10
D19333 N19333 0 diode
R19334 N19333 N19334 10
D19334 N19334 0 diode
R19335 N19334 N19335 10
D19335 N19335 0 diode
R19336 N19335 N19336 10
D19336 N19336 0 diode
R19337 N19336 N19337 10
D19337 N19337 0 diode
R19338 N19337 N19338 10
D19338 N19338 0 diode
R19339 N19338 N19339 10
D19339 N19339 0 diode
R19340 N19339 N19340 10
D19340 N19340 0 diode
R19341 N19340 N19341 10
D19341 N19341 0 diode
R19342 N19341 N19342 10
D19342 N19342 0 diode
R19343 N19342 N19343 10
D19343 N19343 0 diode
R19344 N19343 N19344 10
D19344 N19344 0 diode
R19345 N19344 N19345 10
D19345 N19345 0 diode
R19346 N19345 N19346 10
D19346 N19346 0 diode
R19347 N19346 N19347 10
D19347 N19347 0 diode
R19348 N19347 N19348 10
D19348 N19348 0 diode
R19349 N19348 N19349 10
D19349 N19349 0 diode
R19350 N19349 N19350 10
D19350 N19350 0 diode
R19351 N19350 N19351 10
D19351 N19351 0 diode
R19352 N19351 N19352 10
D19352 N19352 0 diode
R19353 N19352 N19353 10
D19353 N19353 0 diode
R19354 N19353 N19354 10
D19354 N19354 0 diode
R19355 N19354 N19355 10
D19355 N19355 0 diode
R19356 N19355 N19356 10
D19356 N19356 0 diode
R19357 N19356 N19357 10
D19357 N19357 0 diode
R19358 N19357 N19358 10
D19358 N19358 0 diode
R19359 N19358 N19359 10
D19359 N19359 0 diode
R19360 N19359 N19360 10
D19360 N19360 0 diode
R19361 N19360 N19361 10
D19361 N19361 0 diode
R19362 N19361 N19362 10
D19362 N19362 0 diode
R19363 N19362 N19363 10
D19363 N19363 0 diode
R19364 N19363 N19364 10
D19364 N19364 0 diode
R19365 N19364 N19365 10
D19365 N19365 0 diode
R19366 N19365 N19366 10
D19366 N19366 0 diode
R19367 N19366 N19367 10
D19367 N19367 0 diode
R19368 N19367 N19368 10
D19368 N19368 0 diode
R19369 N19368 N19369 10
D19369 N19369 0 diode
R19370 N19369 N19370 10
D19370 N19370 0 diode
R19371 N19370 N19371 10
D19371 N19371 0 diode
R19372 N19371 N19372 10
D19372 N19372 0 diode
R19373 N19372 N19373 10
D19373 N19373 0 diode
R19374 N19373 N19374 10
D19374 N19374 0 diode
R19375 N19374 N19375 10
D19375 N19375 0 diode
R19376 N19375 N19376 10
D19376 N19376 0 diode
R19377 N19376 N19377 10
D19377 N19377 0 diode
R19378 N19377 N19378 10
D19378 N19378 0 diode
R19379 N19378 N19379 10
D19379 N19379 0 diode
R19380 N19379 N19380 10
D19380 N19380 0 diode
R19381 N19380 N19381 10
D19381 N19381 0 diode
R19382 N19381 N19382 10
D19382 N19382 0 diode
R19383 N19382 N19383 10
D19383 N19383 0 diode
R19384 N19383 N19384 10
D19384 N19384 0 diode
R19385 N19384 N19385 10
D19385 N19385 0 diode
R19386 N19385 N19386 10
D19386 N19386 0 diode
R19387 N19386 N19387 10
D19387 N19387 0 diode
R19388 N19387 N19388 10
D19388 N19388 0 diode
R19389 N19388 N19389 10
D19389 N19389 0 diode
R19390 N19389 N19390 10
D19390 N19390 0 diode
R19391 N19390 N19391 10
D19391 N19391 0 diode
R19392 N19391 N19392 10
D19392 N19392 0 diode
R19393 N19392 N19393 10
D19393 N19393 0 diode
R19394 N19393 N19394 10
D19394 N19394 0 diode
R19395 N19394 N19395 10
D19395 N19395 0 diode
R19396 N19395 N19396 10
D19396 N19396 0 diode
R19397 N19396 N19397 10
D19397 N19397 0 diode
R19398 N19397 N19398 10
D19398 N19398 0 diode
R19399 N19398 N19399 10
D19399 N19399 0 diode
R19400 N19399 N19400 10
D19400 N19400 0 diode
R19401 N19400 N19401 10
D19401 N19401 0 diode
R19402 N19401 N19402 10
D19402 N19402 0 diode
R19403 N19402 N19403 10
D19403 N19403 0 diode
R19404 N19403 N19404 10
D19404 N19404 0 diode
R19405 N19404 N19405 10
D19405 N19405 0 diode
R19406 N19405 N19406 10
D19406 N19406 0 diode
R19407 N19406 N19407 10
D19407 N19407 0 diode
R19408 N19407 N19408 10
D19408 N19408 0 diode
R19409 N19408 N19409 10
D19409 N19409 0 diode
R19410 N19409 N19410 10
D19410 N19410 0 diode
R19411 N19410 N19411 10
D19411 N19411 0 diode
R19412 N19411 N19412 10
D19412 N19412 0 diode
R19413 N19412 N19413 10
D19413 N19413 0 diode
R19414 N19413 N19414 10
D19414 N19414 0 diode
R19415 N19414 N19415 10
D19415 N19415 0 diode
R19416 N19415 N19416 10
D19416 N19416 0 diode
R19417 N19416 N19417 10
D19417 N19417 0 diode
R19418 N19417 N19418 10
D19418 N19418 0 diode
R19419 N19418 N19419 10
D19419 N19419 0 diode
R19420 N19419 N19420 10
D19420 N19420 0 diode
R19421 N19420 N19421 10
D19421 N19421 0 diode
R19422 N19421 N19422 10
D19422 N19422 0 diode
R19423 N19422 N19423 10
D19423 N19423 0 diode
R19424 N19423 N19424 10
D19424 N19424 0 diode
R19425 N19424 N19425 10
D19425 N19425 0 diode
R19426 N19425 N19426 10
D19426 N19426 0 diode
R19427 N19426 N19427 10
D19427 N19427 0 diode
R19428 N19427 N19428 10
D19428 N19428 0 diode
R19429 N19428 N19429 10
D19429 N19429 0 diode
R19430 N19429 N19430 10
D19430 N19430 0 diode
R19431 N19430 N19431 10
D19431 N19431 0 diode
R19432 N19431 N19432 10
D19432 N19432 0 diode
R19433 N19432 N19433 10
D19433 N19433 0 diode
R19434 N19433 N19434 10
D19434 N19434 0 diode
R19435 N19434 N19435 10
D19435 N19435 0 diode
R19436 N19435 N19436 10
D19436 N19436 0 diode
R19437 N19436 N19437 10
D19437 N19437 0 diode
R19438 N19437 N19438 10
D19438 N19438 0 diode
R19439 N19438 N19439 10
D19439 N19439 0 diode
R19440 N19439 N19440 10
D19440 N19440 0 diode
R19441 N19440 N19441 10
D19441 N19441 0 diode
R19442 N19441 N19442 10
D19442 N19442 0 diode
R19443 N19442 N19443 10
D19443 N19443 0 diode
R19444 N19443 N19444 10
D19444 N19444 0 diode
R19445 N19444 N19445 10
D19445 N19445 0 diode
R19446 N19445 N19446 10
D19446 N19446 0 diode
R19447 N19446 N19447 10
D19447 N19447 0 diode
R19448 N19447 N19448 10
D19448 N19448 0 diode
R19449 N19448 N19449 10
D19449 N19449 0 diode
R19450 N19449 N19450 10
D19450 N19450 0 diode
R19451 N19450 N19451 10
D19451 N19451 0 diode
R19452 N19451 N19452 10
D19452 N19452 0 diode
R19453 N19452 N19453 10
D19453 N19453 0 diode
R19454 N19453 N19454 10
D19454 N19454 0 diode
R19455 N19454 N19455 10
D19455 N19455 0 diode
R19456 N19455 N19456 10
D19456 N19456 0 diode
R19457 N19456 N19457 10
D19457 N19457 0 diode
R19458 N19457 N19458 10
D19458 N19458 0 diode
R19459 N19458 N19459 10
D19459 N19459 0 diode
R19460 N19459 N19460 10
D19460 N19460 0 diode
R19461 N19460 N19461 10
D19461 N19461 0 diode
R19462 N19461 N19462 10
D19462 N19462 0 diode
R19463 N19462 N19463 10
D19463 N19463 0 diode
R19464 N19463 N19464 10
D19464 N19464 0 diode
R19465 N19464 N19465 10
D19465 N19465 0 diode
R19466 N19465 N19466 10
D19466 N19466 0 diode
R19467 N19466 N19467 10
D19467 N19467 0 diode
R19468 N19467 N19468 10
D19468 N19468 0 diode
R19469 N19468 N19469 10
D19469 N19469 0 diode
R19470 N19469 N19470 10
D19470 N19470 0 diode
R19471 N19470 N19471 10
D19471 N19471 0 diode
R19472 N19471 N19472 10
D19472 N19472 0 diode
R19473 N19472 N19473 10
D19473 N19473 0 diode
R19474 N19473 N19474 10
D19474 N19474 0 diode
R19475 N19474 N19475 10
D19475 N19475 0 diode
R19476 N19475 N19476 10
D19476 N19476 0 diode
R19477 N19476 N19477 10
D19477 N19477 0 diode
R19478 N19477 N19478 10
D19478 N19478 0 diode
R19479 N19478 N19479 10
D19479 N19479 0 diode
R19480 N19479 N19480 10
D19480 N19480 0 diode
R19481 N19480 N19481 10
D19481 N19481 0 diode
R19482 N19481 N19482 10
D19482 N19482 0 diode
R19483 N19482 N19483 10
D19483 N19483 0 diode
R19484 N19483 N19484 10
D19484 N19484 0 diode
R19485 N19484 N19485 10
D19485 N19485 0 diode
R19486 N19485 N19486 10
D19486 N19486 0 diode
R19487 N19486 N19487 10
D19487 N19487 0 diode
R19488 N19487 N19488 10
D19488 N19488 0 diode
R19489 N19488 N19489 10
D19489 N19489 0 diode
R19490 N19489 N19490 10
D19490 N19490 0 diode
R19491 N19490 N19491 10
D19491 N19491 0 diode
R19492 N19491 N19492 10
D19492 N19492 0 diode
R19493 N19492 N19493 10
D19493 N19493 0 diode
R19494 N19493 N19494 10
D19494 N19494 0 diode
R19495 N19494 N19495 10
D19495 N19495 0 diode
R19496 N19495 N19496 10
D19496 N19496 0 diode
R19497 N19496 N19497 10
D19497 N19497 0 diode
R19498 N19497 N19498 10
D19498 N19498 0 diode
R19499 N19498 N19499 10
D19499 N19499 0 diode
R19500 N19499 N19500 10
D19500 N19500 0 diode
R19501 N19500 N19501 10
D19501 N19501 0 diode
R19502 N19501 N19502 10
D19502 N19502 0 diode
R19503 N19502 N19503 10
D19503 N19503 0 diode
R19504 N19503 N19504 10
D19504 N19504 0 diode
R19505 N19504 N19505 10
D19505 N19505 0 diode
R19506 N19505 N19506 10
D19506 N19506 0 diode
R19507 N19506 N19507 10
D19507 N19507 0 diode
R19508 N19507 N19508 10
D19508 N19508 0 diode
R19509 N19508 N19509 10
D19509 N19509 0 diode
R19510 N19509 N19510 10
D19510 N19510 0 diode
R19511 N19510 N19511 10
D19511 N19511 0 diode
R19512 N19511 N19512 10
D19512 N19512 0 diode
R19513 N19512 N19513 10
D19513 N19513 0 diode
R19514 N19513 N19514 10
D19514 N19514 0 diode
R19515 N19514 N19515 10
D19515 N19515 0 diode
R19516 N19515 N19516 10
D19516 N19516 0 diode
R19517 N19516 N19517 10
D19517 N19517 0 diode
R19518 N19517 N19518 10
D19518 N19518 0 diode
R19519 N19518 N19519 10
D19519 N19519 0 diode
R19520 N19519 N19520 10
D19520 N19520 0 diode
R19521 N19520 N19521 10
D19521 N19521 0 diode
R19522 N19521 N19522 10
D19522 N19522 0 diode
R19523 N19522 N19523 10
D19523 N19523 0 diode
R19524 N19523 N19524 10
D19524 N19524 0 diode
R19525 N19524 N19525 10
D19525 N19525 0 diode
R19526 N19525 N19526 10
D19526 N19526 0 diode
R19527 N19526 N19527 10
D19527 N19527 0 diode
R19528 N19527 N19528 10
D19528 N19528 0 diode
R19529 N19528 N19529 10
D19529 N19529 0 diode
R19530 N19529 N19530 10
D19530 N19530 0 diode
R19531 N19530 N19531 10
D19531 N19531 0 diode
R19532 N19531 N19532 10
D19532 N19532 0 diode
R19533 N19532 N19533 10
D19533 N19533 0 diode
R19534 N19533 N19534 10
D19534 N19534 0 diode
R19535 N19534 N19535 10
D19535 N19535 0 diode
R19536 N19535 N19536 10
D19536 N19536 0 diode
R19537 N19536 N19537 10
D19537 N19537 0 diode
R19538 N19537 N19538 10
D19538 N19538 0 diode
R19539 N19538 N19539 10
D19539 N19539 0 diode
R19540 N19539 N19540 10
D19540 N19540 0 diode
R19541 N19540 N19541 10
D19541 N19541 0 diode
R19542 N19541 N19542 10
D19542 N19542 0 diode
R19543 N19542 N19543 10
D19543 N19543 0 diode
R19544 N19543 N19544 10
D19544 N19544 0 diode
R19545 N19544 N19545 10
D19545 N19545 0 diode
R19546 N19545 N19546 10
D19546 N19546 0 diode
R19547 N19546 N19547 10
D19547 N19547 0 diode
R19548 N19547 N19548 10
D19548 N19548 0 diode
R19549 N19548 N19549 10
D19549 N19549 0 diode
R19550 N19549 N19550 10
D19550 N19550 0 diode
R19551 N19550 N19551 10
D19551 N19551 0 diode
R19552 N19551 N19552 10
D19552 N19552 0 diode
R19553 N19552 N19553 10
D19553 N19553 0 diode
R19554 N19553 N19554 10
D19554 N19554 0 diode
R19555 N19554 N19555 10
D19555 N19555 0 diode
R19556 N19555 N19556 10
D19556 N19556 0 diode
R19557 N19556 N19557 10
D19557 N19557 0 diode
R19558 N19557 N19558 10
D19558 N19558 0 diode
R19559 N19558 N19559 10
D19559 N19559 0 diode
R19560 N19559 N19560 10
D19560 N19560 0 diode
R19561 N19560 N19561 10
D19561 N19561 0 diode
R19562 N19561 N19562 10
D19562 N19562 0 diode
R19563 N19562 N19563 10
D19563 N19563 0 diode
R19564 N19563 N19564 10
D19564 N19564 0 diode
R19565 N19564 N19565 10
D19565 N19565 0 diode
R19566 N19565 N19566 10
D19566 N19566 0 diode
R19567 N19566 N19567 10
D19567 N19567 0 diode
R19568 N19567 N19568 10
D19568 N19568 0 diode
R19569 N19568 N19569 10
D19569 N19569 0 diode
R19570 N19569 N19570 10
D19570 N19570 0 diode
R19571 N19570 N19571 10
D19571 N19571 0 diode
R19572 N19571 N19572 10
D19572 N19572 0 diode
R19573 N19572 N19573 10
D19573 N19573 0 diode
R19574 N19573 N19574 10
D19574 N19574 0 diode
R19575 N19574 N19575 10
D19575 N19575 0 diode
R19576 N19575 N19576 10
D19576 N19576 0 diode
R19577 N19576 N19577 10
D19577 N19577 0 diode
R19578 N19577 N19578 10
D19578 N19578 0 diode
R19579 N19578 N19579 10
D19579 N19579 0 diode
R19580 N19579 N19580 10
D19580 N19580 0 diode
R19581 N19580 N19581 10
D19581 N19581 0 diode
R19582 N19581 N19582 10
D19582 N19582 0 diode
R19583 N19582 N19583 10
D19583 N19583 0 diode
R19584 N19583 N19584 10
D19584 N19584 0 diode
R19585 N19584 N19585 10
D19585 N19585 0 diode
R19586 N19585 N19586 10
D19586 N19586 0 diode
R19587 N19586 N19587 10
D19587 N19587 0 diode
R19588 N19587 N19588 10
D19588 N19588 0 diode
R19589 N19588 N19589 10
D19589 N19589 0 diode
R19590 N19589 N19590 10
D19590 N19590 0 diode
R19591 N19590 N19591 10
D19591 N19591 0 diode
R19592 N19591 N19592 10
D19592 N19592 0 diode
R19593 N19592 N19593 10
D19593 N19593 0 diode
R19594 N19593 N19594 10
D19594 N19594 0 diode
R19595 N19594 N19595 10
D19595 N19595 0 diode
R19596 N19595 N19596 10
D19596 N19596 0 diode
R19597 N19596 N19597 10
D19597 N19597 0 diode
R19598 N19597 N19598 10
D19598 N19598 0 diode
R19599 N19598 N19599 10
D19599 N19599 0 diode
R19600 N19599 N19600 10
D19600 N19600 0 diode
R19601 N19600 N19601 10
D19601 N19601 0 diode
R19602 N19601 N19602 10
D19602 N19602 0 diode
R19603 N19602 N19603 10
D19603 N19603 0 diode
R19604 N19603 N19604 10
D19604 N19604 0 diode
R19605 N19604 N19605 10
D19605 N19605 0 diode
R19606 N19605 N19606 10
D19606 N19606 0 diode
R19607 N19606 N19607 10
D19607 N19607 0 diode
R19608 N19607 N19608 10
D19608 N19608 0 diode
R19609 N19608 N19609 10
D19609 N19609 0 diode
R19610 N19609 N19610 10
D19610 N19610 0 diode
R19611 N19610 N19611 10
D19611 N19611 0 diode
R19612 N19611 N19612 10
D19612 N19612 0 diode
R19613 N19612 N19613 10
D19613 N19613 0 diode
R19614 N19613 N19614 10
D19614 N19614 0 diode
R19615 N19614 N19615 10
D19615 N19615 0 diode
R19616 N19615 N19616 10
D19616 N19616 0 diode
R19617 N19616 N19617 10
D19617 N19617 0 diode
R19618 N19617 N19618 10
D19618 N19618 0 diode
R19619 N19618 N19619 10
D19619 N19619 0 diode
R19620 N19619 N19620 10
D19620 N19620 0 diode
R19621 N19620 N19621 10
D19621 N19621 0 diode
R19622 N19621 N19622 10
D19622 N19622 0 diode
R19623 N19622 N19623 10
D19623 N19623 0 diode
R19624 N19623 N19624 10
D19624 N19624 0 diode
R19625 N19624 N19625 10
D19625 N19625 0 diode
R19626 N19625 N19626 10
D19626 N19626 0 diode
R19627 N19626 N19627 10
D19627 N19627 0 diode
R19628 N19627 N19628 10
D19628 N19628 0 diode
R19629 N19628 N19629 10
D19629 N19629 0 diode
R19630 N19629 N19630 10
D19630 N19630 0 diode
R19631 N19630 N19631 10
D19631 N19631 0 diode
R19632 N19631 N19632 10
D19632 N19632 0 diode
R19633 N19632 N19633 10
D19633 N19633 0 diode
R19634 N19633 N19634 10
D19634 N19634 0 diode
R19635 N19634 N19635 10
D19635 N19635 0 diode
R19636 N19635 N19636 10
D19636 N19636 0 diode
R19637 N19636 N19637 10
D19637 N19637 0 diode
R19638 N19637 N19638 10
D19638 N19638 0 diode
R19639 N19638 N19639 10
D19639 N19639 0 diode
R19640 N19639 N19640 10
D19640 N19640 0 diode
R19641 N19640 N19641 10
D19641 N19641 0 diode
R19642 N19641 N19642 10
D19642 N19642 0 diode
R19643 N19642 N19643 10
D19643 N19643 0 diode
R19644 N19643 N19644 10
D19644 N19644 0 diode
R19645 N19644 N19645 10
D19645 N19645 0 diode
R19646 N19645 N19646 10
D19646 N19646 0 diode
R19647 N19646 N19647 10
D19647 N19647 0 diode
R19648 N19647 N19648 10
D19648 N19648 0 diode
R19649 N19648 N19649 10
D19649 N19649 0 diode
R19650 N19649 N19650 10
D19650 N19650 0 diode
R19651 N19650 N19651 10
D19651 N19651 0 diode
R19652 N19651 N19652 10
D19652 N19652 0 diode
R19653 N19652 N19653 10
D19653 N19653 0 diode
R19654 N19653 N19654 10
D19654 N19654 0 diode
R19655 N19654 N19655 10
D19655 N19655 0 diode
R19656 N19655 N19656 10
D19656 N19656 0 diode
R19657 N19656 N19657 10
D19657 N19657 0 diode
R19658 N19657 N19658 10
D19658 N19658 0 diode
R19659 N19658 N19659 10
D19659 N19659 0 diode
R19660 N19659 N19660 10
D19660 N19660 0 diode
R19661 N19660 N19661 10
D19661 N19661 0 diode
R19662 N19661 N19662 10
D19662 N19662 0 diode
R19663 N19662 N19663 10
D19663 N19663 0 diode
R19664 N19663 N19664 10
D19664 N19664 0 diode
R19665 N19664 N19665 10
D19665 N19665 0 diode
R19666 N19665 N19666 10
D19666 N19666 0 diode
R19667 N19666 N19667 10
D19667 N19667 0 diode
R19668 N19667 N19668 10
D19668 N19668 0 diode
R19669 N19668 N19669 10
D19669 N19669 0 diode
R19670 N19669 N19670 10
D19670 N19670 0 diode
R19671 N19670 N19671 10
D19671 N19671 0 diode
R19672 N19671 N19672 10
D19672 N19672 0 diode
R19673 N19672 N19673 10
D19673 N19673 0 diode
R19674 N19673 N19674 10
D19674 N19674 0 diode
R19675 N19674 N19675 10
D19675 N19675 0 diode
R19676 N19675 N19676 10
D19676 N19676 0 diode
R19677 N19676 N19677 10
D19677 N19677 0 diode
R19678 N19677 N19678 10
D19678 N19678 0 diode
R19679 N19678 N19679 10
D19679 N19679 0 diode
R19680 N19679 N19680 10
D19680 N19680 0 diode
R19681 N19680 N19681 10
D19681 N19681 0 diode
R19682 N19681 N19682 10
D19682 N19682 0 diode
R19683 N19682 N19683 10
D19683 N19683 0 diode
R19684 N19683 N19684 10
D19684 N19684 0 diode
R19685 N19684 N19685 10
D19685 N19685 0 diode
R19686 N19685 N19686 10
D19686 N19686 0 diode
R19687 N19686 N19687 10
D19687 N19687 0 diode
R19688 N19687 N19688 10
D19688 N19688 0 diode
R19689 N19688 N19689 10
D19689 N19689 0 diode
R19690 N19689 N19690 10
D19690 N19690 0 diode
R19691 N19690 N19691 10
D19691 N19691 0 diode
R19692 N19691 N19692 10
D19692 N19692 0 diode
R19693 N19692 N19693 10
D19693 N19693 0 diode
R19694 N19693 N19694 10
D19694 N19694 0 diode
R19695 N19694 N19695 10
D19695 N19695 0 diode
R19696 N19695 N19696 10
D19696 N19696 0 diode
R19697 N19696 N19697 10
D19697 N19697 0 diode
R19698 N19697 N19698 10
D19698 N19698 0 diode
R19699 N19698 N19699 10
D19699 N19699 0 diode
R19700 N19699 N19700 10
D19700 N19700 0 diode
R19701 N19700 N19701 10
D19701 N19701 0 diode
R19702 N19701 N19702 10
D19702 N19702 0 diode
R19703 N19702 N19703 10
D19703 N19703 0 diode
R19704 N19703 N19704 10
D19704 N19704 0 diode
R19705 N19704 N19705 10
D19705 N19705 0 diode
R19706 N19705 N19706 10
D19706 N19706 0 diode
R19707 N19706 N19707 10
D19707 N19707 0 diode
R19708 N19707 N19708 10
D19708 N19708 0 diode
R19709 N19708 N19709 10
D19709 N19709 0 diode
R19710 N19709 N19710 10
D19710 N19710 0 diode
R19711 N19710 N19711 10
D19711 N19711 0 diode
R19712 N19711 N19712 10
D19712 N19712 0 diode
R19713 N19712 N19713 10
D19713 N19713 0 diode
R19714 N19713 N19714 10
D19714 N19714 0 diode
R19715 N19714 N19715 10
D19715 N19715 0 diode
R19716 N19715 N19716 10
D19716 N19716 0 diode
R19717 N19716 N19717 10
D19717 N19717 0 diode
R19718 N19717 N19718 10
D19718 N19718 0 diode
R19719 N19718 N19719 10
D19719 N19719 0 diode
R19720 N19719 N19720 10
D19720 N19720 0 diode
R19721 N19720 N19721 10
D19721 N19721 0 diode
R19722 N19721 N19722 10
D19722 N19722 0 diode
R19723 N19722 N19723 10
D19723 N19723 0 diode
R19724 N19723 N19724 10
D19724 N19724 0 diode
R19725 N19724 N19725 10
D19725 N19725 0 diode
R19726 N19725 N19726 10
D19726 N19726 0 diode
R19727 N19726 N19727 10
D19727 N19727 0 diode
R19728 N19727 N19728 10
D19728 N19728 0 diode
R19729 N19728 N19729 10
D19729 N19729 0 diode
R19730 N19729 N19730 10
D19730 N19730 0 diode
R19731 N19730 N19731 10
D19731 N19731 0 diode
R19732 N19731 N19732 10
D19732 N19732 0 diode
R19733 N19732 N19733 10
D19733 N19733 0 diode
R19734 N19733 N19734 10
D19734 N19734 0 diode
R19735 N19734 N19735 10
D19735 N19735 0 diode
R19736 N19735 N19736 10
D19736 N19736 0 diode
R19737 N19736 N19737 10
D19737 N19737 0 diode
R19738 N19737 N19738 10
D19738 N19738 0 diode
R19739 N19738 N19739 10
D19739 N19739 0 diode
R19740 N19739 N19740 10
D19740 N19740 0 diode
R19741 N19740 N19741 10
D19741 N19741 0 diode
R19742 N19741 N19742 10
D19742 N19742 0 diode
R19743 N19742 N19743 10
D19743 N19743 0 diode
R19744 N19743 N19744 10
D19744 N19744 0 diode
R19745 N19744 N19745 10
D19745 N19745 0 diode
R19746 N19745 N19746 10
D19746 N19746 0 diode
R19747 N19746 N19747 10
D19747 N19747 0 diode
R19748 N19747 N19748 10
D19748 N19748 0 diode
R19749 N19748 N19749 10
D19749 N19749 0 diode
R19750 N19749 N19750 10
D19750 N19750 0 diode
R19751 N19750 N19751 10
D19751 N19751 0 diode
R19752 N19751 N19752 10
D19752 N19752 0 diode
R19753 N19752 N19753 10
D19753 N19753 0 diode
R19754 N19753 N19754 10
D19754 N19754 0 diode
R19755 N19754 N19755 10
D19755 N19755 0 diode
R19756 N19755 N19756 10
D19756 N19756 0 diode
R19757 N19756 N19757 10
D19757 N19757 0 diode
R19758 N19757 N19758 10
D19758 N19758 0 diode
R19759 N19758 N19759 10
D19759 N19759 0 diode
R19760 N19759 N19760 10
D19760 N19760 0 diode
R19761 N19760 N19761 10
D19761 N19761 0 diode
R19762 N19761 N19762 10
D19762 N19762 0 diode
R19763 N19762 N19763 10
D19763 N19763 0 diode
R19764 N19763 N19764 10
D19764 N19764 0 diode
R19765 N19764 N19765 10
D19765 N19765 0 diode
R19766 N19765 N19766 10
D19766 N19766 0 diode
R19767 N19766 N19767 10
D19767 N19767 0 diode
R19768 N19767 N19768 10
D19768 N19768 0 diode
R19769 N19768 N19769 10
D19769 N19769 0 diode
R19770 N19769 N19770 10
D19770 N19770 0 diode
R19771 N19770 N19771 10
D19771 N19771 0 diode
R19772 N19771 N19772 10
D19772 N19772 0 diode
R19773 N19772 N19773 10
D19773 N19773 0 diode
R19774 N19773 N19774 10
D19774 N19774 0 diode
R19775 N19774 N19775 10
D19775 N19775 0 diode
R19776 N19775 N19776 10
D19776 N19776 0 diode
R19777 N19776 N19777 10
D19777 N19777 0 diode
R19778 N19777 N19778 10
D19778 N19778 0 diode
R19779 N19778 N19779 10
D19779 N19779 0 diode
R19780 N19779 N19780 10
D19780 N19780 0 diode
R19781 N19780 N19781 10
D19781 N19781 0 diode
R19782 N19781 N19782 10
D19782 N19782 0 diode
R19783 N19782 N19783 10
D19783 N19783 0 diode
R19784 N19783 N19784 10
D19784 N19784 0 diode
R19785 N19784 N19785 10
D19785 N19785 0 diode
R19786 N19785 N19786 10
D19786 N19786 0 diode
R19787 N19786 N19787 10
D19787 N19787 0 diode
R19788 N19787 N19788 10
D19788 N19788 0 diode
R19789 N19788 N19789 10
D19789 N19789 0 diode
R19790 N19789 N19790 10
D19790 N19790 0 diode
R19791 N19790 N19791 10
D19791 N19791 0 diode
R19792 N19791 N19792 10
D19792 N19792 0 diode
R19793 N19792 N19793 10
D19793 N19793 0 diode
R19794 N19793 N19794 10
D19794 N19794 0 diode
R19795 N19794 N19795 10
D19795 N19795 0 diode
R19796 N19795 N19796 10
D19796 N19796 0 diode
R19797 N19796 N19797 10
D19797 N19797 0 diode
R19798 N19797 N19798 10
D19798 N19798 0 diode
R19799 N19798 N19799 10
D19799 N19799 0 diode
R19800 N19799 N19800 10
D19800 N19800 0 diode
R19801 N19800 N19801 10
D19801 N19801 0 diode
R19802 N19801 N19802 10
D19802 N19802 0 diode
R19803 N19802 N19803 10
D19803 N19803 0 diode
R19804 N19803 N19804 10
D19804 N19804 0 diode
R19805 N19804 N19805 10
D19805 N19805 0 diode
R19806 N19805 N19806 10
D19806 N19806 0 diode
R19807 N19806 N19807 10
D19807 N19807 0 diode
R19808 N19807 N19808 10
D19808 N19808 0 diode
R19809 N19808 N19809 10
D19809 N19809 0 diode
R19810 N19809 N19810 10
D19810 N19810 0 diode
R19811 N19810 N19811 10
D19811 N19811 0 diode
R19812 N19811 N19812 10
D19812 N19812 0 diode
R19813 N19812 N19813 10
D19813 N19813 0 diode
R19814 N19813 N19814 10
D19814 N19814 0 diode
R19815 N19814 N19815 10
D19815 N19815 0 diode
R19816 N19815 N19816 10
D19816 N19816 0 diode
R19817 N19816 N19817 10
D19817 N19817 0 diode
R19818 N19817 N19818 10
D19818 N19818 0 diode
R19819 N19818 N19819 10
D19819 N19819 0 diode
R19820 N19819 N19820 10
D19820 N19820 0 diode
R19821 N19820 N19821 10
D19821 N19821 0 diode
R19822 N19821 N19822 10
D19822 N19822 0 diode
R19823 N19822 N19823 10
D19823 N19823 0 diode
R19824 N19823 N19824 10
D19824 N19824 0 diode
R19825 N19824 N19825 10
D19825 N19825 0 diode
R19826 N19825 N19826 10
D19826 N19826 0 diode
R19827 N19826 N19827 10
D19827 N19827 0 diode
R19828 N19827 N19828 10
D19828 N19828 0 diode
R19829 N19828 N19829 10
D19829 N19829 0 diode
R19830 N19829 N19830 10
D19830 N19830 0 diode
R19831 N19830 N19831 10
D19831 N19831 0 diode
R19832 N19831 N19832 10
D19832 N19832 0 diode
R19833 N19832 N19833 10
D19833 N19833 0 diode
R19834 N19833 N19834 10
D19834 N19834 0 diode
R19835 N19834 N19835 10
D19835 N19835 0 diode
R19836 N19835 N19836 10
D19836 N19836 0 diode
R19837 N19836 N19837 10
D19837 N19837 0 diode
R19838 N19837 N19838 10
D19838 N19838 0 diode
R19839 N19838 N19839 10
D19839 N19839 0 diode
R19840 N19839 N19840 10
D19840 N19840 0 diode
R19841 N19840 N19841 10
D19841 N19841 0 diode
R19842 N19841 N19842 10
D19842 N19842 0 diode
R19843 N19842 N19843 10
D19843 N19843 0 diode
R19844 N19843 N19844 10
D19844 N19844 0 diode
R19845 N19844 N19845 10
D19845 N19845 0 diode
R19846 N19845 N19846 10
D19846 N19846 0 diode
R19847 N19846 N19847 10
D19847 N19847 0 diode
R19848 N19847 N19848 10
D19848 N19848 0 diode
R19849 N19848 N19849 10
D19849 N19849 0 diode
R19850 N19849 N19850 10
D19850 N19850 0 diode
R19851 N19850 N19851 10
D19851 N19851 0 diode
R19852 N19851 N19852 10
D19852 N19852 0 diode
R19853 N19852 N19853 10
D19853 N19853 0 diode
R19854 N19853 N19854 10
D19854 N19854 0 diode
R19855 N19854 N19855 10
D19855 N19855 0 diode
R19856 N19855 N19856 10
D19856 N19856 0 diode
R19857 N19856 N19857 10
D19857 N19857 0 diode
R19858 N19857 N19858 10
D19858 N19858 0 diode
R19859 N19858 N19859 10
D19859 N19859 0 diode
R19860 N19859 N19860 10
D19860 N19860 0 diode
R19861 N19860 N19861 10
D19861 N19861 0 diode
R19862 N19861 N19862 10
D19862 N19862 0 diode
R19863 N19862 N19863 10
D19863 N19863 0 diode
R19864 N19863 N19864 10
D19864 N19864 0 diode
R19865 N19864 N19865 10
D19865 N19865 0 diode
R19866 N19865 N19866 10
D19866 N19866 0 diode
R19867 N19866 N19867 10
D19867 N19867 0 diode
R19868 N19867 N19868 10
D19868 N19868 0 diode
R19869 N19868 N19869 10
D19869 N19869 0 diode
R19870 N19869 N19870 10
D19870 N19870 0 diode
R19871 N19870 N19871 10
D19871 N19871 0 diode
R19872 N19871 N19872 10
D19872 N19872 0 diode
R19873 N19872 N19873 10
D19873 N19873 0 diode
R19874 N19873 N19874 10
D19874 N19874 0 diode
R19875 N19874 N19875 10
D19875 N19875 0 diode
R19876 N19875 N19876 10
D19876 N19876 0 diode
R19877 N19876 N19877 10
D19877 N19877 0 diode
R19878 N19877 N19878 10
D19878 N19878 0 diode
R19879 N19878 N19879 10
D19879 N19879 0 diode
R19880 N19879 N19880 10
D19880 N19880 0 diode
R19881 N19880 N19881 10
D19881 N19881 0 diode
R19882 N19881 N19882 10
D19882 N19882 0 diode
R19883 N19882 N19883 10
D19883 N19883 0 diode
R19884 N19883 N19884 10
D19884 N19884 0 diode
R19885 N19884 N19885 10
D19885 N19885 0 diode
R19886 N19885 N19886 10
D19886 N19886 0 diode
R19887 N19886 N19887 10
D19887 N19887 0 diode
R19888 N19887 N19888 10
D19888 N19888 0 diode
R19889 N19888 N19889 10
D19889 N19889 0 diode
R19890 N19889 N19890 10
D19890 N19890 0 diode
R19891 N19890 N19891 10
D19891 N19891 0 diode
R19892 N19891 N19892 10
D19892 N19892 0 diode
R19893 N19892 N19893 10
D19893 N19893 0 diode
R19894 N19893 N19894 10
D19894 N19894 0 diode
R19895 N19894 N19895 10
D19895 N19895 0 diode
R19896 N19895 N19896 10
D19896 N19896 0 diode
R19897 N19896 N19897 10
D19897 N19897 0 diode
R19898 N19897 N19898 10
D19898 N19898 0 diode
R19899 N19898 N19899 10
D19899 N19899 0 diode
R19900 N19899 N19900 10
D19900 N19900 0 diode
R19901 N19900 N19901 10
D19901 N19901 0 diode
R19902 N19901 N19902 10
D19902 N19902 0 diode
R19903 N19902 N19903 10
D19903 N19903 0 diode
R19904 N19903 N19904 10
D19904 N19904 0 diode
R19905 N19904 N19905 10
D19905 N19905 0 diode
R19906 N19905 N19906 10
D19906 N19906 0 diode
R19907 N19906 N19907 10
D19907 N19907 0 diode
R19908 N19907 N19908 10
D19908 N19908 0 diode
R19909 N19908 N19909 10
D19909 N19909 0 diode
R19910 N19909 N19910 10
D19910 N19910 0 diode
R19911 N19910 N19911 10
D19911 N19911 0 diode
R19912 N19911 N19912 10
D19912 N19912 0 diode
R19913 N19912 N19913 10
D19913 N19913 0 diode
R19914 N19913 N19914 10
D19914 N19914 0 diode
R19915 N19914 N19915 10
D19915 N19915 0 diode
R19916 N19915 N19916 10
D19916 N19916 0 diode
R19917 N19916 N19917 10
D19917 N19917 0 diode
R19918 N19917 N19918 10
D19918 N19918 0 diode
R19919 N19918 N19919 10
D19919 N19919 0 diode
R19920 N19919 N19920 10
D19920 N19920 0 diode
R19921 N19920 N19921 10
D19921 N19921 0 diode
R19922 N19921 N19922 10
D19922 N19922 0 diode
R19923 N19922 N19923 10
D19923 N19923 0 diode
R19924 N19923 N19924 10
D19924 N19924 0 diode
R19925 N19924 N19925 10
D19925 N19925 0 diode
R19926 N19925 N19926 10
D19926 N19926 0 diode
R19927 N19926 N19927 10
D19927 N19927 0 diode
R19928 N19927 N19928 10
D19928 N19928 0 diode
R19929 N19928 N19929 10
D19929 N19929 0 diode
R19930 N19929 N19930 10
D19930 N19930 0 diode
R19931 N19930 N19931 10
D19931 N19931 0 diode
R19932 N19931 N19932 10
D19932 N19932 0 diode
R19933 N19932 N19933 10
D19933 N19933 0 diode
R19934 N19933 N19934 10
D19934 N19934 0 diode
R19935 N19934 N19935 10
D19935 N19935 0 diode
R19936 N19935 N19936 10
D19936 N19936 0 diode
R19937 N19936 N19937 10
D19937 N19937 0 diode
R19938 N19937 N19938 10
D19938 N19938 0 diode
R19939 N19938 N19939 10
D19939 N19939 0 diode
R19940 N19939 N19940 10
D19940 N19940 0 diode
R19941 N19940 N19941 10
D19941 N19941 0 diode
R19942 N19941 N19942 10
D19942 N19942 0 diode
R19943 N19942 N19943 10
D19943 N19943 0 diode
R19944 N19943 N19944 10
D19944 N19944 0 diode
R19945 N19944 N19945 10
D19945 N19945 0 diode
R19946 N19945 N19946 10
D19946 N19946 0 diode
R19947 N19946 N19947 10
D19947 N19947 0 diode
R19948 N19947 N19948 10
D19948 N19948 0 diode
R19949 N19948 N19949 10
D19949 N19949 0 diode
R19950 N19949 N19950 10
D19950 N19950 0 diode
R19951 N19950 N19951 10
D19951 N19951 0 diode
R19952 N19951 N19952 10
D19952 N19952 0 diode
R19953 N19952 N19953 10
D19953 N19953 0 diode
R19954 N19953 N19954 10
D19954 N19954 0 diode
R19955 N19954 N19955 10
D19955 N19955 0 diode
R19956 N19955 N19956 10
D19956 N19956 0 diode
R19957 N19956 N19957 10
D19957 N19957 0 diode
R19958 N19957 N19958 10
D19958 N19958 0 diode
R19959 N19958 N19959 10
D19959 N19959 0 diode
R19960 N19959 N19960 10
D19960 N19960 0 diode
R19961 N19960 N19961 10
D19961 N19961 0 diode
R19962 N19961 N19962 10
D19962 N19962 0 diode
R19963 N19962 N19963 10
D19963 N19963 0 diode
R19964 N19963 N19964 10
D19964 N19964 0 diode
R19965 N19964 N19965 10
D19965 N19965 0 diode
R19966 N19965 N19966 10
D19966 N19966 0 diode
R19967 N19966 N19967 10
D19967 N19967 0 diode
R19968 N19967 N19968 10
D19968 N19968 0 diode
R19969 N19968 N19969 10
D19969 N19969 0 diode
R19970 N19969 N19970 10
D19970 N19970 0 diode
R19971 N19970 N19971 10
D19971 N19971 0 diode
R19972 N19971 N19972 10
D19972 N19972 0 diode
R19973 N19972 N19973 10
D19973 N19973 0 diode
R19974 N19973 N19974 10
D19974 N19974 0 diode
R19975 N19974 N19975 10
D19975 N19975 0 diode
R19976 N19975 N19976 10
D19976 N19976 0 diode
R19977 N19976 N19977 10
D19977 N19977 0 diode
R19978 N19977 N19978 10
D19978 N19978 0 diode
R19979 N19978 N19979 10
D19979 N19979 0 diode
R19980 N19979 N19980 10
D19980 N19980 0 diode
R19981 N19980 N19981 10
D19981 N19981 0 diode
R19982 N19981 N19982 10
D19982 N19982 0 diode
R19983 N19982 N19983 10
D19983 N19983 0 diode
R19984 N19983 N19984 10
D19984 N19984 0 diode
R19985 N19984 N19985 10
D19985 N19985 0 diode
R19986 N19985 N19986 10
D19986 N19986 0 diode
R19987 N19986 N19987 10
D19987 N19987 0 diode
R19988 N19987 N19988 10
D19988 N19988 0 diode
R19989 N19988 N19989 10
D19989 N19989 0 diode
R19990 N19989 N19990 10
D19990 N19990 0 diode
R19991 N19990 N19991 10
D19991 N19991 0 diode
R19992 N19991 N19992 10
D19992 N19992 0 diode
R19993 N19992 N19993 10
D19993 N19993 0 diode
R19994 N19993 N19994 10
D19994 N19994 0 diode
R19995 N19994 N19995 10
D19995 N19995 0 diode
R19996 N19995 N19996 10
D19996 N19996 0 diode
R19997 N19996 N19997 10
D19997 N19997 0 diode
R19998 N19997 N19998 10
D19998 N19998 0 diode
R19999 N19998 N19999 10
D19999 N19999 0 diode
R20000 N19999 N20000 10
D20000 N20000 0 diode
R20001 N20000 N20001 10
D20001 N20001 0 diode
R20002 N20001 N20002 10
D20002 N20002 0 diode
R20003 N20002 N20003 10
D20003 N20003 0 diode
R20004 N20003 N20004 10
D20004 N20004 0 diode
R20005 N20004 N20005 10
D20005 N20005 0 diode
R20006 N20005 N20006 10
D20006 N20006 0 diode
R20007 N20006 N20007 10
D20007 N20007 0 diode
R20008 N20007 N20008 10
D20008 N20008 0 diode
R20009 N20008 N20009 10
D20009 N20009 0 diode
R20010 N20009 N20010 10
D20010 N20010 0 diode
R20011 N20010 N20011 10
D20011 N20011 0 diode
R20012 N20011 N20012 10
D20012 N20012 0 diode
R20013 N20012 N20013 10
D20013 N20013 0 diode
R20014 N20013 N20014 10
D20014 N20014 0 diode
R20015 N20014 N20015 10
D20015 N20015 0 diode
R20016 N20015 N20016 10
D20016 N20016 0 diode
R20017 N20016 N20017 10
D20017 N20017 0 diode
R20018 N20017 N20018 10
D20018 N20018 0 diode
R20019 N20018 N20019 10
D20019 N20019 0 diode
R20020 N20019 N20020 10
D20020 N20020 0 diode
R20021 N20020 N20021 10
D20021 N20021 0 diode
R20022 N20021 N20022 10
D20022 N20022 0 diode
R20023 N20022 N20023 10
D20023 N20023 0 diode
R20024 N20023 N20024 10
D20024 N20024 0 diode
R20025 N20024 N20025 10
D20025 N20025 0 diode
R20026 N20025 N20026 10
D20026 N20026 0 diode
R20027 N20026 N20027 10
D20027 N20027 0 diode
R20028 N20027 N20028 10
D20028 N20028 0 diode
R20029 N20028 N20029 10
D20029 N20029 0 diode
R20030 N20029 N20030 10
D20030 N20030 0 diode
R20031 N20030 N20031 10
D20031 N20031 0 diode
R20032 N20031 N20032 10
D20032 N20032 0 diode
R20033 N20032 N20033 10
D20033 N20033 0 diode
R20034 N20033 N20034 10
D20034 N20034 0 diode
R20035 N20034 N20035 10
D20035 N20035 0 diode
R20036 N20035 N20036 10
D20036 N20036 0 diode
R20037 N20036 N20037 10
D20037 N20037 0 diode
R20038 N20037 N20038 10
D20038 N20038 0 diode
R20039 N20038 N20039 10
D20039 N20039 0 diode
R20040 N20039 N20040 10
D20040 N20040 0 diode
R20041 N20040 N20041 10
D20041 N20041 0 diode
R20042 N20041 N20042 10
D20042 N20042 0 diode
R20043 N20042 N20043 10
D20043 N20043 0 diode
R20044 N20043 N20044 10
D20044 N20044 0 diode
R20045 N20044 N20045 10
D20045 N20045 0 diode
R20046 N20045 N20046 10
D20046 N20046 0 diode
R20047 N20046 N20047 10
D20047 N20047 0 diode
R20048 N20047 N20048 10
D20048 N20048 0 diode
R20049 N20048 N20049 10
D20049 N20049 0 diode
R20050 N20049 N20050 10
D20050 N20050 0 diode
R20051 N20050 N20051 10
D20051 N20051 0 diode
R20052 N20051 N20052 10
D20052 N20052 0 diode
R20053 N20052 N20053 10
D20053 N20053 0 diode
R20054 N20053 N20054 10
D20054 N20054 0 diode
R20055 N20054 N20055 10
D20055 N20055 0 diode
R20056 N20055 N20056 10
D20056 N20056 0 diode
R20057 N20056 N20057 10
D20057 N20057 0 diode
R20058 N20057 N20058 10
D20058 N20058 0 diode
R20059 N20058 N20059 10
D20059 N20059 0 diode
R20060 N20059 N20060 10
D20060 N20060 0 diode
R20061 N20060 N20061 10
D20061 N20061 0 diode
R20062 N20061 N20062 10
D20062 N20062 0 diode
R20063 N20062 N20063 10
D20063 N20063 0 diode
R20064 N20063 N20064 10
D20064 N20064 0 diode
R20065 N20064 N20065 10
D20065 N20065 0 diode
R20066 N20065 N20066 10
D20066 N20066 0 diode
R20067 N20066 N20067 10
D20067 N20067 0 diode
R20068 N20067 N20068 10
D20068 N20068 0 diode
R20069 N20068 N20069 10
D20069 N20069 0 diode
R20070 N20069 N20070 10
D20070 N20070 0 diode
R20071 N20070 N20071 10
D20071 N20071 0 diode
R20072 N20071 N20072 10
D20072 N20072 0 diode
R20073 N20072 N20073 10
D20073 N20073 0 diode
R20074 N20073 N20074 10
D20074 N20074 0 diode
R20075 N20074 N20075 10
D20075 N20075 0 diode
R20076 N20075 N20076 10
D20076 N20076 0 diode
R20077 N20076 N20077 10
D20077 N20077 0 diode
R20078 N20077 N20078 10
D20078 N20078 0 diode
R20079 N20078 N20079 10
D20079 N20079 0 diode
R20080 N20079 N20080 10
D20080 N20080 0 diode
R20081 N20080 N20081 10
D20081 N20081 0 diode
R20082 N20081 N20082 10
D20082 N20082 0 diode
R20083 N20082 N20083 10
D20083 N20083 0 diode
R20084 N20083 N20084 10
D20084 N20084 0 diode
R20085 N20084 N20085 10
D20085 N20085 0 diode
R20086 N20085 N20086 10
D20086 N20086 0 diode
R20087 N20086 N20087 10
D20087 N20087 0 diode
R20088 N20087 N20088 10
D20088 N20088 0 diode
R20089 N20088 N20089 10
D20089 N20089 0 diode
R20090 N20089 N20090 10
D20090 N20090 0 diode
R20091 N20090 N20091 10
D20091 N20091 0 diode
R20092 N20091 N20092 10
D20092 N20092 0 diode
R20093 N20092 N20093 10
D20093 N20093 0 diode
R20094 N20093 N20094 10
D20094 N20094 0 diode
R20095 N20094 N20095 10
D20095 N20095 0 diode
R20096 N20095 N20096 10
D20096 N20096 0 diode
R20097 N20096 N20097 10
D20097 N20097 0 diode
R20098 N20097 N20098 10
D20098 N20098 0 diode
R20099 N20098 N20099 10
D20099 N20099 0 diode
R20100 N20099 N20100 10
D20100 N20100 0 diode
R20101 N20100 N20101 10
D20101 N20101 0 diode
R20102 N20101 N20102 10
D20102 N20102 0 diode
R20103 N20102 N20103 10
D20103 N20103 0 diode
R20104 N20103 N20104 10
D20104 N20104 0 diode
R20105 N20104 N20105 10
D20105 N20105 0 diode
R20106 N20105 N20106 10
D20106 N20106 0 diode
R20107 N20106 N20107 10
D20107 N20107 0 diode
R20108 N20107 N20108 10
D20108 N20108 0 diode
R20109 N20108 N20109 10
D20109 N20109 0 diode
R20110 N20109 N20110 10
D20110 N20110 0 diode
R20111 N20110 N20111 10
D20111 N20111 0 diode
R20112 N20111 N20112 10
D20112 N20112 0 diode
R20113 N20112 N20113 10
D20113 N20113 0 diode
R20114 N20113 N20114 10
D20114 N20114 0 diode
R20115 N20114 N20115 10
D20115 N20115 0 diode
R20116 N20115 N20116 10
D20116 N20116 0 diode
R20117 N20116 N20117 10
D20117 N20117 0 diode
R20118 N20117 N20118 10
D20118 N20118 0 diode
R20119 N20118 N20119 10
D20119 N20119 0 diode
R20120 N20119 N20120 10
D20120 N20120 0 diode
R20121 N20120 N20121 10
D20121 N20121 0 diode
R20122 N20121 N20122 10
D20122 N20122 0 diode
R20123 N20122 N20123 10
D20123 N20123 0 diode
R20124 N20123 N20124 10
D20124 N20124 0 diode
R20125 N20124 N20125 10
D20125 N20125 0 diode
R20126 N20125 N20126 10
D20126 N20126 0 diode
R20127 N20126 N20127 10
D20127 N20127 0 diode
R20128 N20127 N20128 10
D20128 N20128 0 diode
R20129 N20128 N20129 10
D20129 N20129 0 diode
R20130 N20129 N20130 10
D20130 N20130 0 diode
R20131 N20130 N20131 10
D20131 N20131 0 diode
R20132 N20131 N20132 10
D20132 N20132 0 diode
R20133 N20132 N20133 10
D20133 N20133 0 diode
R20134 N20133 N20134 10
D20134 N20134 0 diode
R20135 N20134 N20135 10
D20135 N20135 0 diode
R20136 N20135 N20136 10
D20136 N20136 0 diode
R20137 N20136 N20137 10
D20137 N20137 0 diode
R20138 N20137 N20138 10
D20138 N20138 0 diode
R20139 N20138 N20139 10
D20139 N20139 0 diode
R20140 N20139 N20140 10
D20140 N20140 0 diode
R20141 N20140 N20141 10
D20141 N20141 0 diode
R20142 N20141 N20142 10
D20142 N20142 0 diode
R20143 N20142 N20143 10
D20143 N20143 0 diode
R20144 N20143 N20144 10
D20144 N20144 0 diode
R20145 N20144 N20145 10
D20145 N20145 0 diode
R20146 N20145 N20146 10
D20146 N20146 0 diode
R20147 N20146 N20147 10
D20147 N20147 0 diode
R20148 N20147 N20148 10
D20148 N20148 0 diode
R20149 N20148 N20149 10
D20149 N20149 0 diode
R20150 N20149 N20150 10
D20150 N20150 0 diode
R20151 N20150 N20151 10
D20151 N20151 0 diode
R20152 N20151 N20152 10
D20152 N20152 0 diode
R20153 N20152 N20153 10
D20153 N20153 0 diode
R20154 N20153 N20154 10
D20154 N20154 0 diode
R20155 N20154 N20155 10
D20155 N20155 0 diode
R20156 N20155 N20156 10
D20156 N20156 0 diode
R20157 N20156 N20157 10
D20157 N20157 0 diode
R20158 N20157 N20158 10
D20158 N20158 0 diode
R20159 N20158 N20159 10
D20159 N20159 0 diode
R20160 N20159 N20160 10
D20160 N20160 0 diode
R20161 N20160 N20161 10
D20161 N20161 0 diode
R20162 N20161 N20162 10
D20162 N20162 0 diode
R20163 N20162 N20163 10
D20163 N20163 0 diode
R20164 N20163 N20164 10
D20164 N20164 0 diode
R20165 N20164 N20165 10
D20165 N20165 0 diode
R20166 N20165 N20166 10
D20166 N20166 0 diode
R20167 N20166 N20167 10
D20167 N20167 0 diode
R20168 N20167 N20168 10
D20168 N20168 0 diode
R20169 N20168 N20169 10
D20169 N20169 0 diode
R20170 N20169 N20170 10
D20170 N20170 0 diode
R20171 N20170 N20171 10
D20171 N20171 0 diode
R20172 N20171 N20172 10
D20172 N20172 0 diode
R20173 N20172 N20173 10
D20173 N20173 0 diode
R20174 N20173 N20174 10
D20174 N20174 0 diode
R20175 N20174 N20175 10
D20175 N20175 0 diode
R20176 N20175 N20176 10
D20176 N20176 0 diode
R20177 N20176 N20177 10
D20177 N20177 0 diode
R20178 N20177 N20178 10
D20178 N20178 0 diode
R20179 N20178 N20179 10
D20179 N20179 0 diode
R20180 N20179 N20180 10
D20180 N20180 0 diode
R20181 N20180 N20181 10
D20181 N20181 0 diode
R20182 N20181 N20182 10
D20182 N20182 0 diode
R20183 N20182 N20183 10
D20183 N20183 0 diode
R20184 N20183 N20184 10
D20184 N20184 0 diode
R20185 N20184 N20185 10
D20185 N20185 0 diode
R20186 N20185 N20186 10
D20186 N20186 0 diode
R20187 N20186 N20187 10
D20187 N20187 0 diode
R20188 N20187 N20188 10
D20188 N20188 0 diode
R20189 N20188 N20189 10
D20189 N20189 0 diode
R20190 N20189 N20190 10
D20190 N20190 0 diode
R20191 N20190 N20191 10
D20191 N20191 0 diode
R20192 N20191 N20192 10
D20192 N20192 0 diode
R20193 N20192 N20193 10
D20193 N20193 0 diode
R20194 N20193 N20194 10
D20194 N20194 0 diode
R20195 N20194 N20195 10
D20195 N20195 0 diode
R20196 N20195 N20196 10
D20196 N20196 0 diode
R20197 N20196 N20197 10
D20197 N20197 0 diode
R20198 N20197 N20198 10
D20198 N20198 0 diode
R20199 N20198 N20199 10
D20199 N20199 0 diode
R20200 N20199 N20200 10
D20200 N20200 0 diode
R20201 N20200 N20201 10
D20201 N20201 0 diode
R20202 N20201 N20202 10
D20202 N20202 0 diode
R20203 N20202 N20203 10
D20203 N20203 0 diode
R20204 N20203 N20204 10
D20204 N20204 0 diode
R20205 N20204 N20205 10
D20205 N20205 0 diode
R20206 N20205 N20206 10
D20206 N20206 0 diode
R20207 N20206 N20207 10
D20207 N20207 0 diode
R20208 N20207 N20208 10
D20208 N20208 0 diode
R20209 N20208 N20209 10
D20209 N20209 0 diode
R20210 N20209 N20210 10
D20210 N20210 0 diode
R20211 N20210 N20211 10
D20211 N20211 0 diode
R20212 N20211 N20212 10
D20212 N20212 0 diode
R20213 N20212 N20213 10
D20213 N20213 0 diode
R20214 N20213 N20214 10
D20214 N20214 0 diode
R20215 N20214 N20215 10
D20215 N20215 0 diode
R20216 N20215 N20216 10
D20216 N20216 0 diode
R20217 N20216 N20217 10
D20217 N20217 0 diode
R20218 N20217 N20218 10
D20218 N20218 0 diode
R20219 N20218 N20219 10
D20219 N20219 0 diode
R20220 N20219 N20220 10
D20220 N20220 0 diode
R20221 N20220 N20221 10
D20221 N20221 0 diode
R20222 N20221 N20222 10
D20222 N20222 0 diode
R20223 N20222 N20223 10
D20223 N20223 0 diode
R20224 N20223 N20224 10
D20224 N20224 0 diode
R20225 N20224 N20225 10
D20225 N20225 0 diode
R20226 N20225 N20226 10
D20226 N20226 0 diode
R20227 N20226 N20227 10
D20227 N20227 0 diode
R20228 N20227 N20228 10
D20228 N20228 0 diode
R20229 N20228 N20229 10
D20229 N20229 0 diode
R20230 N20229 N20230 10
D20230 N20230 0 diode
R20231 N20230 N20231 10
D20231 N20231 0 diode
R20232 N20231 N20232 10
D20232 N20232 0 diode
R20233 N20232 N20233 10
D20233 N20233 0 diode
R20234 N20233 N20234 10
D20234 N20234 0 diode
R20235 N20234 N20235 10
D20235 N20235 0 diode
R20236 N20235 N20236 10
D20236 N20236 0 diode
R20237 N20236 N20237 10
D20237 N20237 0 diode
R20238 N20237 N20238 10
D20238 N20238 0 diode
R20239 N20238 N20239 10
D20239 N20239 0 diode
R20240 N20239 N20240 10
D20240 N20240 0 diode
R20241 N20240 N20241 10
D20241 N20241 0 diode
R20242 N20241 N20242 10
D20242 N20242 0 diode
R20243 N20242 N20243 10
D20243 N20243 0 diode
R20244 N20243 N20244 10
D20244 N20244 0 diode
R20245 N20244 N20245 10
D20245 N20245 0 diode
R20246 N20245 N20246 10
D20246 N20246 0 diode
R20247 N20246 N20247 10
D20247 N20247 0 diode
R20248 N20247 N20248 10
D20248 N20248 0 diode
R20249 N20248 N20249 10
D20249 N20249 0 diode
R20250 N20249 N20250 10
D20250 N20250 0 diode
R20251 N20250 N20251 10
D20251 N20251 0 diode
R20252 N20251 N20252 10
D20252 N20252 0 diode
R20253 N20252 N20253 10
D20253 N20253 0 diode
R20254 N20253 N20254 10
D20254 N20254 0 diode
R20255 N20254 N20255 10
D20255 N20255 0 diode
R20256 N20255 N20256 10
D20256 N20256 0 diode
R20257 N20256 N20257 10
D20257 N20257 0 diode
R20258 N20257 N20258 10
D20258 N20258 0 diode
R20259 N20258 N20259 10
D20259 N20259 0 diode
R20260 N20259 N20260 10
D20260 N20260 0 diode
R20261 N20260 N20261 10
D20261 N20261 0 diode
R20262 N20261 N20262 10
D20262 N20262 0 diode
R20263 N20262 N20263 10
D20263 N20263 0 diode
R20264 N20263 N20264 10
D20264 N20264 0 diode
R20265 N20264 N20265 10
D20265 N20265 0 diode
R20266 N20265 N20266 10
D20266 N20266 0 diode
R20267 N20266 N20267 10
D20267 N20267 0 diode
R20268 N20267 N20268 10
D20268 N20268 0 diode
R20269 N20268 N20269 10
D20269 N20269 0 diode
R20270 N20269 N20270 10
D20270 N20270 0 diode
R20271 N20270 N20271 10
D20271 N20271 0 diode
R20272 N20271 N20272 10
D20272 N20272 0 diode
R20273 N20272 N20273 10
D20273 N20273 0 diode
R20274 N20273 N20274 10
D20274 N20274 0 diode
R20275 N20274 N20275 10
D20275 N20275 0 diode
R20276 N20275 N20276 10
D20276 N20276 0 diode
R20277 N20276 N20277 10
D20277 N20277 0 diode
R20278 N20277 N20278 10
D20278 N20278 0 diode
R20279 N20278 N20279 10
D20279 N20279 0 diode
R20280 N20279 N20280 10
D20280 N20280 0 diode
R20281 N20280 N20281 10
D20281 N20281 0 diode
R20282 N20281 N20282 10
D20282 N20282 0 diode
R20283 N20282 N20283 10
D20283 N20283 0 diode
R20284 N20283 N20284 10
D20284 N20284 0 diode
R20285 N20284 N20285 10
D20285 N20285 0 diode
R20286 N20285 N20286 10
D20286 N20286 0 diode
R20287 N20286 N20287 10
D20287 N20287 0 diode
R20288 N20287 N20288 10
D20288 N20288 0 diode
R20289 N20288 N20289 10
D20289 N20289 0 diode
R20290 N20289 N20290 10
D20290 N20290 0 diode
R20291 N20290 N20291 10
D20291 N20291 0 diode
R20292 N20291 N20292 10
D20292 N20292 0 diode
R20293 N20292 N20293 10
D20293 N20293 0 diode
R20294 N20293 N20294 10
D20294 N20294 0 diode
R20295 N20294 N20295 10
D20295 N20295 0 diode
R20296 N20295 N20296 10
D20296 N20296 0 diode
R20297 N20296 N20297 10
D20297 N20297 0 diode
R20298 N20297 N20298 10
D20298 N20298 0 diode
R20299 N20298 N20299 10
D20299 N20299 0 diode
R20300 N20299 N20300 10
D20300 N20300 0 diode
R20301 N20300 N20301 10
D20301 N20301 0 diode
R20302 N20301 N20302 10
D20302 N20302 0 diode
R20303 N20302 N20303 10
D20303 N20303 0 diode
R20304 N20303 N20304 10
D20304 N20304 0 diode
R20305 N20304 N20305 10
D20305 N20305 0 diode
R20306 N20305 N20306 10
D20306 N20306 0 diode
R20307 N20306 N20307 10
D20307 N20307 0 diode
R20308 N20307 N20308 10
D20308 N20308 0 diode
R20309 N20308 N20309 10
D20309 N20309 0 diode
R20310 N20309 N20310 10
D20310 N20310 0 diode
R20311 N20310 N20311 10
D20311 N20311 0 diode
R20312 N20311 N20312 10
D20312 N20312 0 diode
R20313 N20312 N20313 10
D20313 N20313 0 diode
R20314 N20313 N20314 10
D20314 N20314 0 diode
R20315 N20314 N20315 10
D20315 N20315 0 diode
R20316 N20315 N20316 10
D20316 N20316 0 diode
R20317 N20316 N20317 10
D20317 N20317 0 diode
R20318 N20317 N20318 10
D20318 N20318 0 diode
R20319 N20318 N20319 10
D20319 N20319 0 diode
R20320 N20319 N20320 10
D20320 N20320 0 diode
R20321 N20320 N20321 10
D20321 N20321 0 diode
R20322 N20321 N20322 10
D20322 N20322 0 diode
R20323 N20322 N20323 10
D20323 N20323 0 diode
R20324 N20323 N20324 10
D20324 N20324 0 diode
R20325 N20324 N20325 10
D20325 N20325 0 diode
R20326 N20325 N20326 10
D20326 N20326 0 diode
R20327 N20326 N20327 10
D20327 N20327 0 diode
R20328 N20327 N20328 10
D20328 N20328 0 diode
R20329 N20328 N20329 10
D20329 N20329 0 diode
R20330 N20329 N20330 10
D20330 N20330 0 diode
R20331 N20330 N20331 10
D20331 N20331 0 diode
R20332 N20331 N20332 10
D20332 N20332 0 diode
R20333 N20332 N20333 10
D20333 N20333 0 diode
R20334 N20333 N20334 10
D20334 N20334 0 diode
R20335 N20334 N20335 10
D20335 N20335 0 diode
R20336 N20335 N20336 10
D20336 N20336 0 diode
R20337 N20336 N20337 10
D20337 N20337 0 diode
R20338 N20337 N20338 10
D20338 N20338 0 diode
R20339 N20338 N20339 10
D20339 N20339 0 diode
R20340 N20339 N20340 10
D20340 N20340 0 diode
R20341 N20340 N20341 10
D20341 N20341 0 diode
R20342 N20341 N20342 10
D20342 N20342 0 diode
R20343 N20342 N20343 10
D20343 N20343 0 diode
R20344 N20343 N20344 10
D20344 N20344 0 diode
R20345 N20344 N20345 10
D20345 N20345 0 diode
R20346 N20345 N20346 10
D20346 N20346 0 diode
R20347 N20346 N20347 10
D20347 N20347 0 diode
R20348 N20347 N20348 10
D20348 N20348 0 diode
R20349 N20348 N20349 10
D20349 N20349 0 diode
R20350 N20349 N20350 10
D20350 N20350 0 diode
R20351 N20350 N20351 10
D20351 N20351 0 diode
R20352 N20351 N20352 10
D20352 N20352 0 diode
R20353 N20352 N20353 10
D20353 N20353 0 diode
R20354 N20353 N20354 10
D20354 N20354 0 diode
R20355 N20354 N20355 10
D20355 N20355 0 diode
R20356 N20355 N20356 10
D20356 N20356 0 diode
R20357 N20356 N20357 10
D20357 N20357 0 diode
R20358 N20357 N20358 10
D20358 N20358 0 diode
R20359 N20358 N20359 10
D20359 N20359 0 diode
R20360 N20359 N20360 10
D20360 N20360 0 diode
R20361 N20360 N20361 10
D20361 N20361 0 diode
R20362 N20361 N20362 10
D20362 N20362 0 diode
R20363 N20362 N20363 10
D20363 N20363 0 diode
R20364 N20363 N20364 10
D20364 N20364 0 diode
R20365 N20364 N20365 10
D20365 N20365 0 diode
R20366 N20365 N20366 10
D20366 N20366 0 diode
R20367 N20366 N20367 10
D20367 N20367 0 diode
R20368 N20367 N20368 10
D20368 N20368 0 diode
R20369 N20368 N20369 10
D20369 N20369 0 diode
R20370 N20369 N20370 10
D20370 N20370 0 diode
R20371 N20370 N20371 10
D20371 N20371 0 diode
R20372 N20371 N20372 10
D20372 N20372 0 diode
R20373 N20372 N20373 10
D20373 N20373 0 diode
R20374 N20373 N20374 10
D20374 N20374 0 diode
R20375 N20374 N20375 10
D20375 N20375 0 diode
R20376 N20375 N20376 10
D20376 N20376 0 diode
R20377 N20376 N20377 10
D20377 N20377 0 diode
R20378 N20377 N20378 10
D20378 N20378 0 diode
R20379 N20378 N20379 10
D20379 N20379 0 diode
R20380 N20379 N20380 10
D20380 N20380 0 diode
R20381 N20380 N20381 10
D20381 N20381 0 diode
R20382 N20381 N20382 10
D20382 N20382 0 diode
R20383 N20382 N20383 10
D20383 N20383 0 diode
R20384 N20383 N20384 10
D20384 N20384 0 diode
R20385 N20384 N20385 10
D20385 N20385 0 diode
R20386 N20385 N20386 10
D20386 N20386 0 diode
R20387 N20386 N20387 10
D20387 N20387 0 diode
R20388 N20387 N20388 10
D20388 N20388 0 diode
R20389 N20388 N20389 10
D20389 N20389 0 diode
R20390 N20389 N20390 10
D20390 N20390 0 diode
R20391 N20390 N20391 10
D20391 N20391 0 diode
R20392 N20391 N20392 10
D20392 N20392 0 diode
R20393 N20392 N20393 10
D20393 N20393 0 diode
R20394 N20393 N20394 10
D20394 N20394 0 diode
R20395 N20394 N20395 10
D20395 N20395 0 diode
R20396 N20395 N20396 10
D20396 N20396 0 diode
R20397 N20396 N20397 10
D20397 N20397 0 diode
R20398 N20397 N20398 10
D20398 N20398 0 diode
R20399 N20398 N20399 10
D20399 N20399 0 diode
R20400 N20399 N20400 10
D20400 N20400 0 diode
R20401 N20400 N20401 10
D20401 N20401 0 diode
R20402 N20401 N20402 10
D20402 N20402 0 diode
R20403 N20402 N20403 10
D20403 N20403 0 diode
R20404 N20403 N20404 10
D20404 N20404 0 diode
R20405 N20404 N20405 10
D20405 N20405 0 diode
R20406 N20405 N20406 10
D20406 N20406 0 diode
R20407 N20406 N20407 10
D20407 N20407 0 diode
R20408 N20407 N20408 10
D20408 N20408 0 diode
R20409 N20408 N20409 10
D20409 N20409 0 diode
R20410 N20409 N20410 10
D20410 N20410 0 diode
R20411 N20410 N20411 10
D20411 N20411 0 diode
R20412 N20411 N20412 10
D20412 N20412 0 diode
R20413 N20412 N20413 10
D20413 N20413 0 diode
R20414 N20413 N20414 10
D20414 N20414 0 diode
R20415 N20414 N20415 10
D20415 N20415 0 diode
R20416 N20415 N20416 10
D20416 N20416 0 diode
R20417 N20416 N20417 10
D20417 N20417 0 diode
R20418 N20417 N20418 10
D20418 N20418 0 diode
R20419 N20418 N20419 10
D20419 N20419 0 diode
R20420 N20419 N20420 10
D20420 N20420 0 diode
R20421 N20420 N20421 10
D20421 N20421 0 diode
R20422 N20421 N20422 10
D20422 N20422 0 diode
R20423 N20422 N20423 10
D20423 N20423 0 diode
R20424 N20423 N20424 10
D20424 N20424 0 diode
R20425 N20424 N20425 10
D20425 N20425 0 diode
R20426 N20425 N20426 10
D20426 N20426 0 diode
R20427 N20426 N20427 10
D20427 N20427 0 diode
R20428 N20427 N20428 10
D20428 N20428 0 diode
R20429 N20428 N20429 10
D20429 N20429 0 diode
R20430 N20429 N20430 10
D20430 N20430 0 diode
R20431 N20430 N20431 10
D20431 N20431 0 diode
R20432 N20431 N20432 10
D20432 N20432 0 diode
R20433 N20432 N20433 10
D20433 N20433 0 diode
R20434 N20433 N20434 10
D20434 N20434 0 diode
R20435 N20434 N20435 10
D20435 N20435 0 diode
R20436 N20435 N20436 10
D20436 N20436 0 diode
R20437 N20436 N20437 10
D20437 N20437 0 diode
R20438 N20437 N20438 10
D20438 N20438 0 diode
R20439 N20438 N20439 10
D20439 N20439 0 diode
R20440 N20439 N20440 10
D20440 N20440 0 diode
R20441 N20440 N20441 10
D20441 N20441 0 diode
R20442 N20441 N20442 10
D20442 N20442 0 diode
R20443 N20442 N20443 10
D20443 N20443 0 diode
R20444 N20443 N20444 10
D20444 N20444 0 diode
R20445 N20444 N20445 10
D20445 N20445 0 diode
R20446 N20445 N20446 10
D20446 N20446 0 diode
R20447 N20446 N20447 10
D20447 N20447 0 diode
R20448 N20447 N20448 10
D20448 N20448 0 diode
R20449 N20448 N20449 10
D20449 N20449 0 diode
R20450 N20449 N20450 10
D20450 N20450 0 diode
R20451 N20450 N20451 10
D20451 N20451 0 diode
R20452 N20451 N20452 10
D20452 N20452 0 diode
R20453 N20452 N20453 10
D20453 N20453 0 diode
R20454 N20453 N20454 10
D20454 N20454 0 diode
R20455 N20454 N20455 10
D20455 N20455 0 diode
R20456 N20455 N20456 10
D20456 N20456 0 diode
R20457 N20456 N20457 10
D20457 N20457 0 diode
R20458 N20457 N20458 10
D20458 N20458 0 diode
R20459 N20458 N20459 10
D20459 N20459 0 diode
R20460 N20459 N20460 10
D20460 N20460 0 diode
R20461 N20460 N20461 10
D20461 N20461 0 diode
R20462 N20461 N20462 10
D20462 N20462 0 diode
R20463 N20462 N20463 10
D20463 N20463 0 diode
R20464 N20463 N20464 10
D20464 N20464 0 diode
R20465 N20464 N20465 10
D20465 N20465 0 diode
R20466 N20465 N20466 10
D20466 N20466 0 diode
R20467 N20466 N20467 10
D20467 N20467 0 diode
R20468 N20467 N20468 10
D20468 N20468 0 diode
R20469 N20468 N20469 10
D20469 N20469 0 diode
R20470 N20469 N20470 10
D20470 N20470 0 diode
R20471 N20470 N20471 10
D20471 N20471 0 diode
R20472 N20471 N20472 10
D20472 N20472 0 diode
R20473 N20472 N20473 10
D20473 N20473 0 diode
R20474 N20473 N20474 10
D20474 N20474 0 diode
R20475 N20474 N20475 10
D20475 N20475 0 diode
R20476 N20475 N20476 10
D20476 N20476 0 diode
R20477 N20476 N20477 10
D20477 N20477 0 diode
R20478 N20477 N20478 10
D20478 N20478 0 diode
R20479 N20478 N20479 10
D20479 N20479 0 diode
R20480 N20479 N20480 10
D20480 N20480 0 diode
R20481 N20480 N20481 10
D20481 N20481 0 diode
R20482 N20481 N20482 10
D20482 N20482 0 diode
R20483 N20482 N20483 10
D20483 N20483 0 diode
R20484 N20483 N20484 10
D20484 N20484 0 diode
R20485 N20484 N20485 10
D20485 N20485 0 diode
R20486 N20485 N20486 10
D20486 N20486 0 diode
R20487 N20486 N20487 10
D20487 N20487 0 diode
R20488 N20487 N20488 10
D20488 N20488 0 diode
R20489 N20488 N20489 10
D20489 N20489 0 diode
R20490 N20489 N20490 10
D20490 N20490 0 diode
R20491 N20490 N20491 10
D20491 N20491 0 diode
R20492 N20491 N20492 10
D20492 N20492 0 diode
R20493 N20492 N20493 10
D20493 N20493 0 diode
R20494 N20493 N20494 10
D20494 N20494 0 diode
R20495 N20494 N20495 10
D20495 N20495 0 diode
R20496 N20495 N20496 10
D20496 N20496 0 diode
R20497 N20496 N20497 10
D20497 N20497 0 diode
R20498 N20497 N20498 10
D20498 N20498 0 diode
R20499 N20498 N20499 10
D20499 N20499 0 diode
R20500 N20499 N20500 10
D20500 N20500 0 diode
R20501 N20500 N20501 10
D20501 N20501 0 diode
R20502 N20501 N20502 10
D20502 N20502 0 diode
R20503 N20502 N20503 10
D20503 N20503 0 diode
R20504 N20503 N20504 10
D20504 N20504 0 diode
R20505 N20504 N20505 10
D20505 N20505 0 diode
R20506 N20505 N20506 10
D20506 N20506 0 diode
R20507 N20506 N20507 10
D20507 N20507 0 diode
R20508 N20507 N20508 10
D20508 N20508 0 diode
R20509 N20508 N20509 10
D20509 N20509 0 diode
R20510 N20509 N20510 10
D20510 N20510 0 diode
R20511 N20510 N20511 10
D20511 N20511 0 diode
R20512 N20511 N20512 10
D20512 N20512 0 diode
R20513 N20512 N20513 10
D20513 N20513 0 diode
R20514 N20513 N20514 10
D20514 N20514 0 diode
R20515 N20514 N20515 10
D20515 N20515 0 diode
R20516 N20515 N20516 10
D20516 N20516 0 diode
R20517 N20516 N20517 10
D20517 N20517 0 diode
R20518 N20517 N20518 10
D20518 N20518 0 diode
R20519 N20518 N20519 10
D20519 N20519 0 diode
R20520 N20519 N20520 10
D20520 N20520 0 diode
R20521 N20520 N20521 10
D20521 N20521 0 diode
R20522 N20521 N20522 10
D20522 N20522 0 diode
R20523 N20522 N20523 10
D20523 N20523 0 diode
R20524 N20523 N20524 10
D20524 N20524 0 diode
R20525 N20524 N20525 10
D20525 N20525 0 diode
R20526 N20525 N20526 10
D20526 N20526 0 diode
R20527 N20526 N20527 10
D20527 N20527 0 diode
R20528 N20527 N20528 10
D20528 N20528 0 diode
R20529 N20528 N20529 10
D20529 N20529 0 diode
R20530 N20529 N20530 10
D20530 N20530 0 diode
R20531 N20530 N20531 10
D20531 N20531 0 diode
R20532 N20531 N20532 10
D20532 N20532 0 diode
R20533 N20532 N20533 10
D20533 N20533 0 diode
R20534 N20533 N20534 10
D20534 N20534 0 diode
R20535 N20534 N20535 10
D20535 N20535 0 diode
R20536 N20535 N20536 10
D20536 N20536 0 diode
R20537 N20536 N20537 10
D20537 N20537 0 diode
R20538 N20537 N20538 10
D20538 N20538 0 diode
R20539 N20538 N20539 10
D20539 N20539 0 diode
R20540 N20539 N20540 10
D20540 N20540 0 diode
R20541 N20540 N20541 10
D20541 N20541 0 diode
R20542 N20541 N20542 10
D20542 N20542 0 diode
R20543 N20542 N20543 10
D20543 N20543 0 diode
R20544 N20543 N20544 10
D20544 N20544 0 diode
R20545 N20544 N20545 10
D20545 N20545 0 diode
R20546 N20545 N20546 10
D20546 N20546 0 diode
R20547 N20546 N20547 10
D20547 N20547 0 diode
R20548 N20547 N20548 10
D20548 N20548 0 diode
R20549 N20548 N20549 10
D20549 N20549 0 diode
R20550 N20549 N20550 10
D20550 N20550 0 diode
R20551 N20550 N20551 10
D20551 N20551 0 diode
R20552 N20551 N20552 10
D20552 N20552 0 diode
R20553 N20552 N20553 10
D20553 N20553 0 diode
R20554 N20553 N20554 10
D20554 N20554 0 diode
R20555 N20554 N20555 10
D20555 N20555 0 diode
R20556 N20555 N20556 10
D20556 N20556 0 diode
R20557 N20556 N20557 10
D20557 N20557 0 diode
R20558 N20557 N20558 10
D20558 N20558 0 diode
R20559 N20558 N20559 10
D20559 N20559 0 diode
R20560 N20559 N20560 10
D20560 N20560 0 diode
R20561 N20560 N20561 10
D20561 N20561 0 diode
R20562 N20561 N20562 10
D20562 N20562 0 diode
R20563 N20562 N20563 10
D20563 N20563 0 diode
R20564 N20563 N20564 10
D20564 N20564 0 diode
R20565 N20564 N20565 10
D20565 N20565 0 diode
R20566 N20565 N20566 10
D20566 N20566 0 diode
R20567 N20566 N20567 10
D20567 N20567 0 diode
R20568 N20567 N20568 10
D20568 N20568 0 diode
R20569 N20568 N20569 10
D20569 N20569 0 diode
R20570 N20569 N20570 10
D20570 N20570 0 diode
R20571 N20570 N20571 10
D20571 N20571 0 diode
R20572 N20571 N20572 10
D20572 N20572 0 diode
R20573 N20572 N20573 10
D20573 N20573 0 diode
R20574 N20573 N20574 10
D20574 N20574 0 diode
R20575 N20574 N20575 10
D20575 N20575 0 diode
R20576 N20575 N20576 10
D20576 N20576 0 diode
R20577 N20576 N20577 10
D20577 N20577 0 diode
R20578 N20577 N20578 10
D20578 N20578 0 diode
R20579 N20578 N20579 10
D20579 N20579 0 diode
R20580 N20579 N20580 10
D20580 N20580 0 diode
R20581 N20580 N20581 10
D20581 N20581 0 diode
R20582 N20581 N20582 10
D20582 N20582 0 diode
R20583 N20582 N20583 10
D20583 N20583 0 diode
R20584 N20583 N20584 10
D20584 N20584 0 diode
R20585 N20584 N20585 10
D20585 N20585 0 diode
R20586 N20585 N20586 10
D20586 N20586 0 diode
R20587 N20586 N20587 10
D20587 N20587 0 diode
R20588 N20587 N20588 10
D20588 N20588 0 diode
R20589 N20588 N20589 10
D20589 N20589 0 diode
R20590 N20589 N20590 10
D20590 N20590 0 diode
R20591 N20590 N20591 10
D20591 N20591 0 diode
R20592 N20591 N20592 10
D20592 N20592 0 diode
R20593 N20592 N20593 10
D20593 N20593 0 diode
R20594 N20593 N20594 10
D20594 N20594 0 diode
R20595 N20594 N20595 10
D20595 N20595 0 diode
R20596 N20595 N20596 10
D20596 N20596 0 diode
R20597 N20596 N20597 10
D20597 N20597 0 diode
R20598 N20597 N20598 10
D20598 N20598 0 diode
R20599 N20598 N20599 10
D20599 N20599 0 diode
R20600 N20599 N20600 10
D20600 N20600 0 diode
R20601 N20600 N20601 10
D20601 N20601 0 diode
R20602 N20601 N20602 10
D20602 N20602 0 diode
R20603 N20602 N20603 10
D20603 N20603 0 diode
R20604 N20603 N20604 10
D20604 N20604 0 diode
R20605 N20604 N20605 10
D20605 N20605 0 diode
R20606 N20605 N20606 10
D20606 N20606 0 diode
R20607 N20606 N20607 10
D20607 N20607 0 diode
R20608 N20607 N20608 10
D20608 N20608 0 diode
R20609 N20608 N20609 10
D20609 N20609 0 diode
R20610 N20609 N20610 10
D20610 N20610 0 diode
R20611 N20610 N20611 10
D20611 N20611 0 diode
R20612 N20611 N20612 10
D20612 N20612 0 diode
R20613 N20612 N20613 10
D20613 N20613 0 diode
R20614 N20613 N20614 10
D20614 N20614 0 diode
R20615 N20614 N20615 10
D20615 N20615 0 diode
R20616 N20615 N20616 10
D20616 N20616 0 diode
R20617 N20616 N20617 10
D20617 N20617 0 diode
R20618 N20617 N20618 10
D20618 N20618 0 diode
R20619 N20618 N20619 10
D20619 N20619 0 diode
R20620 N20619 N20620 10
D20620 N20620 0 diode
R20621 N20620 N20621 10
D20621 N20621 0 diode
R20622 N20621 N20622 10
D20622 N20622 0 diode
R20623 N20622 N20623 10
D20623 N20623 0 diode
R20624 N20623 N20624 10
D20624 N20624 0 diode
R20625 N20624 N20625 10
D20625 N20625 0 diode
R20626 N20625 N20626 10
D20626 N20626 0 diode
R20627 N20626 N20627 10
D20627 N20627 0 diode
R20628 N20627 N20628 10
D20628 N20628 0 diode
R20629 N20628 N20629 10
D20629 N20629 0 diode
R20630 N20629 N20630 10
D20630 N20630 0 diode
R20631 N20630 N20631 10
D20631 N20631 0 diode
R20632 N20631 N20632 10
D20632 N20632 0 diode
R20633 N20632 N20633 10
D20633 N20633 0 diode
R20634 N20633 N20634 10
D20634 N20634 0 diode
R20635 N20634 N20635 10
D20635 N20635 0 diode
R20636 N20635 N20636 10
D20636 N20636 0 diode
R20637 N20636 N20637 10
D20637 N20637 0 diode
R20638 N20637 N20638 10
D20638 N20638 0 diode
R20639 N20638 N20639 10
D20639 N20639 0 diode
R20640 N20639 N20640 10
D20640 N20640 0 diode
R20641 N20640 N20641 10
D20641 N20641 0 diode
R20642 N20641 N20642 10
D20642 N20642 0 diode
R20643 N20642 N20643 10
D20643 N20643 0 diode
R20644 N20643 N20644 10
D20644 N20644 0 diode
R20645 N20644 N20645 10
D20645 N20645 0 diode
R20646 N20645 N20646 10
D20646 N20646 0 diode
R20647 N20646 N20647 10
D20647 N20647 0 diode
R20648 N20647 N20648 10
D20648 N20648 0 diode
R20649 N20648 N20649 10
D20649 N20649 0 diode
R20650 N20649 N20650 10
D20650 N20650 0 diode
R20651 N20650 N20651 10
D20651 N20651 0 diode
R20652 N20651 N20652 10
D20652 N20652 0 diode
R20653 N20652 N20653 10
D20653 N20653 0 diode
R20654 N20653 N20654 10
D20654 N20654 0 diode
R20655 N20654 N20655 10
D20655 N20655 0 diode
R20656 N20655 N20656 10
D20656 N20656 0 diode
R20657 N20656 N20657 10
D20657 N20657 0 diode
R20658 N20657 N20658 10
D20658 N20658 0 diode
R20659 N20658 N20659 10
D20659 N20659 0 diode
R20660 N20659 N20660 10
D20660 N20660 0 diode
R20661 N20660 N20661 10
D20661 N20661 0 diode
R20662 N20661 N20662 10
D20662 N20662 0 diode
R20663 N20662 N20663 10
D20663 N20663 0 diode
R20664 N20663 N20664 10
D20664 N20664 0 diode
R20665 N20664 N20665 10
D20665 N20665 0 diode
R20666 N20665 N20666 10
D20666 N20666 0 diode
R20667 N20666 N20667 10
D20667 N20667 0 diode
R20668 N20667 N20668 10
D20668 N20668 0 diode
R20669 N20668 N20669 10
D20669 N20669 0 diode
R20670 N20669 N20670 10
D20670 N20670 0 diode
R20671 N20670 N20671 10
D20671 N20671 0 diode
R20672 N20671 N20672 10
D20672 N20672 0 diode
R20673 N20672 N20673 10
D20673 N20673 0 diode
R20674 N20673 N20674 10
D20674 N20674 0 diode
R20675 N20674 N20675 10
D20675 N20675 0 diode
R20676 N20675 N20676 10
D20676 N20676 0 diode
R20677 N20676 N20677 10
D20677 N20677 0 diode
R20678 N20677 N20678 10
D20678 N20678 0 diode
R20679 N20678 N20679 10
D20679 N20679 0 diode
R20680 N20679 N20680 10
D20680 N20680 0 diode
R20681 N20680 N20681 10
D20681 N20681 0 diode
R20682 N20681 N20682 10
D20682 N20682 0 diode
R20683 N20682 N20683 10
D20683 N20683 0 diode
R20684 N20683 N20684 10
D20684 N20684 0 diode
R20685 N20684 N20685 10
D20685 N20685 0 diode
R20686 N20685 N20686 10
D20686 N20686 0 diode
R20687 N20686 N20687 10
D20687 N20687 0 diode
R20688 N20687 N20688 10
D20688 N20688 0 diode
R20689 N20688 N20689 10
D20689 N20689 0 diode
R20690 N20689 N20690 10
D20690 N20690 0 diode
R20691 N20690 N20691 10
D20691 N20691 0 diode
R20692 N20691 N20692 10
D20692 N20692 0 diode
R20693 N20692 N20693 10
D20693 N20693 0 diode
R20694 N20693 N20694 10
D20694 N20694 0 diode
R20695 N20694 N20695 10
D20695 N20695 0 diode
R20696 N20695 N20696 10
D20696 N20696 0 diode
R20697 N20696 N20697 10
D20697 N20697 0 diode
R20698 N20697 N20698 10
D20698 N20698 0 diode
R20699 N20698 N20699 10
D20699 N20699 0 diode
R20700 N20699 N20700 10
D20700 N20700 0 diode
R20701 N20700 N20701 10
D20701 N20701 0 diode
R20702 N20701 N20702 10
D20702 N20702 0 diode
R20703 N20702 N20703 10
D20703 N20703 0 diode
R20704 N20703 N20704 10
D20704 N20704 0 diode
R20705 N20704 N20705 10
D20705 N20705 0 diode
R20706 N20705 N20706 10
D20706 N20706 0 diode
R20707 N20706 N20707 10
D20707 N20707 0 diode
R20708 N20707 N20708 10
D20708 N20708 0 diode
R20709 N20708 N20709 10
D20709 N20709 0 diode
R20710 N20709 N20710 10
D20710 N20710 0 diode
R20711 N20710 N20711 10
D20711 N20711 0 diode
R20712 N20711 N20712 10
D20712 N20712 0 diode
R20713 N20712 N20713 10
D20713 N20713 0 diode
R20714 N20713 N20714 10
D20714 N20714 0 diode
R20715 N20714 N20715 10
D20715 N20715 0 diode
R20716 N20715 N20716 10
D20716 N20716 0 diode
R20717 N20716 N20717 10
D20717 N20717 0 diode
R20718 N20717 N20718 10
D20718 N20718 0 diode
R20719 N20718 N20719 10
D20719 N20719 0 diode
R20720 N20719 N20720 10
D20720 N20720 0 diode
R20721 N20720 N20721 10
D20721 N20721 0 diode
R20722 N20721 N20722 10
D20722 N20722 0 diode
R20723 N20722 N20723 10
D20723 N20723 0 diode
R20724 N20723 N20724 10
D20724 N20724 0 diode
R20725 N20724 N20725 10
D20725 N20725 0 diode
R20726 N20725 N20726 10
D20726 N20726 0 diode
R20727 N20726 N20727 10
D20727 N20727 0 diode
R20728 N20727 N20728 10
D20728 N20728 0 diode
R20729 N20728 N20729 10
D20729 N20729 0 diode
R20730 N20729 N20730 10
D20730 N20730 0 diode
R20731 N20730 N20731 10
D20731 N20731 0 diode
R20732 N20731 N20732 10
D20732 N20732 0 diode
R20733 N20732 N20733 10
D20733 N20733 0 diode
R20734 N20733 N20734 10
D20734 N20734 0 diode
R20735 N20734 N20735 10
D20735 N20735 0 diode
R20736 N20735 N20736 10
D20736 N20736 0 diode
R20737 N20736 N20737 10
D20737 N20737 0 diode
R20738 N20737 N20738 10
D20738 N20738 0 diode
R20739 N20738 N20739 10
D20739 N20739 0 diode
R20740 N20739 N20740 10
D20740 N20740 0 diode
R20741 N20740 N20741 10
D20741 N20741 0 diode
R20742 N20741 N20742 10
D20742 N20742 0 diode
R20743 N20742 N20743 10
D20743 N20743 0 diode
R20744 N20743 N20744 10
D20744 N20744 0 diode
R20745 N20744 N20745 10
D20745 N20745 0 diode
R20746 N20745 N20746 10
D20746 N20746 0 diode
R20747 N20746 N20747 10
D20747 N20747 0 diode
R20748 N20747 N20748 10
D20748 N20748 0 diode
R20749 N20748 N20749 10
D20749 N20749 0 diode
R20750 N20749 N20750 10
D20750 N20750 0 diode
R20751 N20750 N20751 10
D20751 N20751 0 diode
R20752 N20751 N20752 10
D20752 N20752 0 diode
R20753 N20752 N20753 10
D20753 N20753 0 diode
R20754 N20753 N20754 10
D20754 N20754 0 diode
R20755 N20754 N20755 10
D20755 N20755 0 diode
R20756 N20755 N20756 10
D20756 N20756 0 diode
R20757 N20756 N20757 10
D20757 N20757 0 diode
R20758 N20757 N20758 10
D20758 N20758 0 diode
R20759 N20758 N20759 10
D20759 N20759 0 diode
R20760 N20759 N20760 10
D20760 N20760 0 diode
R20761 N20760 N20761 10
D20761 N20761 0 diode
R20762 N20761 N20762 10
D20762 N20762 0 diode
R20763 N20762 N20763 10
D20763 N20763 0 diode
R20764 N20763 N20764 10
D20764 N20764 0 diode
R20765 N20764 N20765 10
D20765 N20765 0 diode
R20766 N20765 N20766 10
D20766 N20766 0 diode
R20767 N20766 N20767 10
D20767 N20767 0 diode
R20768 N20767 N20768 10
D20768 N20768 0 diode
R20769 N20768 N20769 10
D20769 N20769 0 diode
R20770 N20769 N20770 10
D20770 N20770 0 diode
R20771 N20770 N20771 10
D20771 N20771 0 diode
R20772 N20771 N20772 10
D20772 N20772 0 diode
R20773 N20772 N20773 10
D20773 N20773 0 diode
R20774 N20773 N20774 10
D20774 N20774 0 diode
R20775 N20774 N20775 10
D20775 N20775 0 diode
R20776 N20775 N20776 10
D20776 N20776 0 diode
R20777 N20776 N20777 10
D20777 N20777 0 diode
R20778 N20777 N20778 10
D20778 N20778 0 diode
R20779 N20778 N20779 10
D20779 N20779 0 diode
R20780 N20779 N20780 10
D20780 N20780 0 diode
R20781 N20780 N20781 10
D20781 N20781 0 diode
R20782 N20781 N20782 10
D20782 N20782 0 diode
R20783 N20782 N20783 10
D20783 N20783 0 diode
R20784 N20783 N20784 10
D20784 N20784 0 diode
R20785 N20784 N20785 10
D20785 N20785 0 diode
R20786 N20785 N20786 10
D20786 N20786 0 diode
R20787 N20786 N20787 10
D20787 N20787 0 diode
R20788 N20787 N20788 10
D20788 N20788 0 diode
R20789 N20788 N20789 10
D20789 N20789 0 diode
R20790 N20789 N20790 10
D20790 N20790 0 diode
R20791 N20790 N20791 10
D20791 N20791 0 diode
R20792 N20791 N20792 10
D20792 N20792 0 diode
R20793 N20792 N20793 10
D20793 N20793 0 diode
R20794 N20793 N20794 10
D20794 N20794 0 diode
R20795 N20794 N20795 10
D20795 N20795 0 diode
R20796 N20795 N20796 10
D20796 N20796 0 diode
R20797 N20796 N20797 10
D20797 N20797 0 diode
R20798 N20797 N20798 10
D20798 N20798 0 diode
R20799 N20798 N20799 10
D20799 N20799 0 diode
R20800 N20799 N20800 10
D20800 N20800 0 diode
R20801 N20800 N20801 10
D20801 N20801 0 diode
R20802 N20801 N20802 10
D20802 N20802 0 diode
R20803 N20802 N20803 10
D20803 N20803 0 diode
R20804 N20803 N20804 10
D20804 N20804 0 diode
R20805 N20804 N20805 10
D20805 N20805 0 diode
R20806 N20805 N20806 10
D20806 N20806 0 diode
R20807 N20806 N20807 10
D20807 N20807 0 diode
R20808 N20807 N20808 10
D20808 N20808 0 diode
R20809 N20808 N20809 10
D20809 N20809 0 diode
R20810 N20809 N20810 10
D20810 N20810 0 diode
R20811 N20810 N20811 10
D20811 N20811 0 diode
R20812 N20811 N20812 10
D20812 N20812 0 diode
R20813 N20812 N20813 10
D20813 N20813 0 diode
R20814 N20813 N20814 10
D20814 N20814 0 diode
R20815 N20814 N20815 10
D20815 N20815 0 diode
R20816 N20815 N20816 10
D20816 N20816 0 diode
R20817 N20816 N20817 10
D20817 N20817 0 diode
R20818 N20817 N20818 10
D20818 N20818 0 diode
R20819 N20818 N20819 10
D20819 N20819 0 diode
R20820 N20819 N20820 10
D20820 N20820 0 diode
R20821 N20820 N20821 10
D20821 N20821 0 diode
R20822 N20821 N20822 10
D20822 N20822 0 diode
R20823 N20822 N20823 10
D20823 N20823 0 diode
R20824 N20823 N20824 10
D20824 N20824 0 diode
R20825 N20824 N20825 10
D20825 N20825 0 diode
R20826 N20825 N20826 10
D20826 N20826 0 diode
R20827 N20826 N20827 10
D20827 N20827 0 diode
R20828 N20827 N20828 10
D20828 N20828 0 diode
R20829 N20828 N20829 10
D20829 N20829 0 diode
R20830 N20829 N20830 10
D20830 N20830 0 diode
R20831 N20830 N20831 10
D20831 N20831 0 diode
R20832 N20831 N20832 10
D20832 N20832 0 diode
R20833 N20832 N20833 10
D20833 N20833 0 diode
R20834 N20833 N20834 10
D20834 N20834 0 diode
R20835 N20834 N20835 10
D20835 N20835 0 diode
R20836 N20835 N20836 10
D20836 N20836 0 diode
R20837 N20836 N20837 10
D20837 N20837 0 diode
R20838 N20837 N20838 10
D20838 N20838 0 diode
R20839 N20838 N20839 10
D20839 N20839 0 diode
R20840 N20839 N20840 10
D20840 N20840 0 diode
R20841 N20840 N20841 10
D20841 N20841 0 diode
R20842 N20841 N20842 10
D20842 N20842 0 diode
R20843 N20842 N20843 10
D20843 N20843 0 diode
R20844 N20843 N20844 10
D20844 N20844 0 diode
R20845 N20844 N20845 10
D20845 N20845 0 diode
R20846 N20845 N20846 10
D20846 N20846 0 diode
R20847 N20846 N20847 10
D20847 N20847 0 diode
R20848 N20847 N20848 10
D20848 N20848 0 diode
R20849 N20848 N20849 10
D20849 N20849 0 diode
R20850 N20849 N20850 10
D20850 N20850 0 diode
R20851 N20850 N20851 10
D20851 N20851 0 diode
R20852 N20851 N20852 10
D20852 N20852 0 diode
R20853 N20852 N20853 10
D20853 N20853 0 diode
R20854 N20853 N20854 10
D20854 N20854 0 diode
R20855 N20854 N20855 10
D20855 N20855 0 diode
R20856 N20855 N20856 10
D20856 N20856 0 diode
R20857 N20856 N20857 10
D20857 N20857 0 diode
R20858 N20857 N20858 10
D20858 N20858 0 diode
R20859 N20858 N20859 10
D20859 N20859 0 diode
R20860 N20859 N20860 10
D20860 N20860 0 diode
R20861 N20860 N20861 10
D20861 N20861 0 diode
R20862 N20861 N20862 10
D20862 N20862 0 diode
R20863 N20862 N20863 10
D20863 N20863 0 diode
R20864 N20863 N20864 10
D20864 N20864 0 diode
R20865 N20864 N20865 10
D20865 N20865 0 diode
R20866 N20865 N20866 10
D20866 N20866 0 diode
R20867 N20866 N20867 10
D20867 N20867 0 diode
R20868 N20867 N20868 10
D20868 N20868 0 diode
R20869 N20868 N20869 10
D20869 N20869 0 diode
R20870 N20869 N20870 10
D20870 N20870 0 diode
R20871 N20870 N20871 10
D20871 N20871 0 diode
R20872 N20871 N20872 10
D20872 N20872 0 diode
R20873 N20872 N20873 10
D20873 N20873 0 diode
R20874 N20873 N20874 10
D20874 N20874 0 diode
R20875 N20874 N20875 10
D20875 N20875 0 diode
R20876 N20875 N20876 10
D20876 N20876 0 diode
R20877 N20876 N20877 10
D20877 N20877 0 diode
R20878 N20877 N20878 10
D20878 N20878 0 diode
R20879 N20878 N20879 10
D20879 N20879 0 diode
R20880 N20879 N20880 10
D20880 N20880 0 diode
R20881 N20880 N20881 10
D20881 N20881 0 diode
R20882 N20881 N20882 10
D20882 N20882 0 diode
R20883 N20882 N20883 10
D20883 N20883 0 diode
R20884 N20883 N20884 10
D20884 N20884 0 diode
R20885 N20884 N20885 10
D20885 N20885 0 diode
R20886 N20885 N20886 10
D20886 N20886 0 diode
R20887 N20886 N20887 10
D20887 N20887 0 diode
R20888 N20887 N20888 10
D20888 N20888 0 diode
R20889 N20888 N20889 10
D20889 N20889 0 diode
R20890 N20889 N20890 10
D20890 N20890 0 diode
R20891 N20890 N20891 10
D20891 N20891 0 diode
R20892 N20891 N20892 10
D20892 N20892 0 diode
R20893 N20892 N20893 10
D20893 N20893 0 diode
R20894 N20893 N20894 10
D20894 N20894 0 diode
R20895 N20894 N20895 10
D20895 N20895 0 diode
R20896 N20895 N20896 10
D20896 N20896 0 diode
R20897 N20896 N20897 10
D20897 N20897 0 diode
R20898 N20897 N20898 10
D20898 N20898 0 diode
R20899 N20898 N20899 10
D20899 N20899 0 diode
R20900 N20899 N20900 10
D20900 N20900 0 diode
R20901 N20900 N20901 10
D20901 N20901 0 diode
R20902 N20901 N20902 10
D20902 N20902 0 diode
R20903 N20902 N20903 10
D20903 N20903 0 diode
R20904 N20903 N20904 10
D20904 N20904 0 diode
R20905 N20904 N20905 10
D20905 N20905 0 diode
R20906 N20905 N20906 10
D20906 N20906 0 diode
R20907 N20906 N20907 10
D20907 N20907 0 diode
R20908 N20907 N20908 10
D20908 N20908 0 diode
R20909 N20908 N20909 10
D20909 N20909 0 diode
R20910 N20909 N20910 10
D20910 N20910 0 diode
R20911 N20910 N20911 10
D20911 N20911 0 diode
R20912 N20911 N20912 10
D20912 N20912 0 diode
R20913 N20912 N20913 10
D20913 N20913 0 diode
R20914 N20913 N20914 10
D20914 N20914 0 diode
R20915 N20914 N20915 10
D20915 N20915 0 diode
R20916 N20915 N20916 10
D20916 N20916 0 diode
R20917 N20916 N20917 10
D20917 N20917 0 diode
R20918 N20917 N20918 10
D20918 N20918 0 diode
R20919 N20918 N20919 10
D20919 N20919 0 diode
R20920 N20919 N20920 10
D20920 N20920 0 diode
R20921 N20920 N20921 10
D20921 N20921 0 diode
R20922 N20921 N20922 10
D20922 N20922 0 diode
R20923 N20922 N20923 10
D20923 N20923 0 diode
R20924 N20923 N20924 10
D20924 N20924 0 diode
R20925 N20924 N20925 10
D20925 N20925 0 diode
R20926 N20925 N20926 10
D20926 N20926 0 diode
R20927 N20926 N20927 10
D20927 N20927 0 diode
R20928 N20927 N20928 10
D20928 N20928 0 diode
R20929 N20928 N20929 10
D20929 N20929 0 diode
R20930 N20929 N20930 10
D20930 N20930 0 diode
R20931 N20930 N20931 10
D20931 N20931 0 diode
R20932 N20931 N20932 10
D20932 N20932 0 diode
R20933 N20932 N20933 10
D20933 N20933 0 diode
R20934 N20933 N20934 10
D20934 N20934 0 diode
R20935 N20934 N20935 10
D20935 N20935 0 diode
R20936 N20935 N20936 10
D20936 N20936 0 diode
R20937 N20936 N20937 10
D20937 N20937 0 diode
R20938 N20937 N20938 10
D20938 N20938 0 diode
R20939 N20938 N20939 10
D20939 N20939 0 diode
R20940 N20939 N20940 10
D20940 N20940 0 diode
R20941 N20940 N20941 10
D20941 N20941 0 diode
R20942 N20941 N20942 10
D20942 N20942 0 diode
R20943 N20942 N20943 10
D20943 N20943 0 diode
R20944 N20943 N20944 10
D20944 N20944 0 diode
R20945 N20944 N20945 10
D20945 N20945 0 diode
R20946 N20945 N20946 10
D20946 N20946 0 diode
R20947 N20946 N20947 10
D20947 N20947 0 diode
R20948 N20947 N20948 10
D20948 N20948 0 diode
R20949 N20948 N20949 10
D20949 N20949 0 diode
R20950 N20949 N20950 10
D20950 N20950 0 diode
R20951 N20950 N20951 10
D20951 N20951 0 diode
R20952 N20951 N20952 10
D20952 N20952 0 diode
R20953 N20952 N20953 10
D20953 N20953 0 diode
R20954 N20953 N20954 10
D20954 N20954 0 diode
R20955 N20954 N20955 10
D20955 N20955 0 diode
R20956 N20955 N20956 10
D20956 N20956 0 diode
R20957 N20956 N20957 10
D20957 N20957 0 diode
R20958 N20957 N20958 10
D20958 N20958 0 diode
R20959 N20958 N20959 10
D20959 N20959 0 diode
R20960 N20959 N20960 10
D20960 N20960 0 diode
R20961 N20960 N20961 10
D20961 N20961 0 diode
R20962 N20961 N20962 10
D20962 N20962 0 diode
R20963 N20962 N20963 10
D20963 N20963 0 diode
R20964 N20963 N20964 10
D20964 N20964 0 diode
R20965 N20964 N20965 10
D20965 N20965 0 diode
R20966 N20965 N20966 10
D20966 N20966 0 diode
R20967 N20966 N20967 10
D20967 N20967 0 diode
R20968 N20967 N20968 10
D20968 N20968 0 diode
R20969 N20968 N20969 10
D20969 N20969 0 diode
R20970 N20969 N20970 10
D20970 N20970 0 diode
R20971 N20970 N20971 10
D20971 N20971 0 diode
R20972 N20971 N20972 10
D20972 N20972 0 diode
R20973 N20972 N20973 10
D20973 N20973 0 diode
R20974 N20973 N20974 10
D20974 N20974 0 diode
R20975 N20974 N20975 10
D20975 N20975 0 diode
R20976 N20975 N20976 10
D20976 N20976 0 diode
R20977 N20976 N20977 10
D20977 N20977 0 diode
R20978 N20977 N20978 10
D20978 N20978 0 diode
R20979 N20978 N20979 10
D20979 N20979 0 diode
R20980 N20979 N20980 10
D20980 N20980 0 diode
R20981 N20980 N20981 10
D20981 N20981 0 diode
R20982 N20981 N20982 10
D20982 N20982 0 diode
R20983 N20982 N20983 10
D20983 N20983 0 diode
R20984 N20983 N20984 10
D20984 N20984 0 diode
R20985 N20984 N20985 10
D20985 N20985 0 diode
R20986 N20985 N20986 10
D20986 N20986 0 diode
R20987 N20986 N20987 10
D20987 N20987 0 diode
R20988 N20987 N20988 10
D20988 N20988 0 diode
R20989 N20988 N20989 10
D20989 N20989 0 diode
R20990 N20989 N20990 10
D20990 N20990 0 diode
R20991 N20990 N20991 10
D20991 N20991 0 diode
R20992 N20991 N20992 10
D20992 N20992 0 diode
R20993 N20992 N20993 10
D20993 N20993 0 diode
R20994 N20993 N20994 10
D20994 N20994 0 diode
R20995 N20994 N20995 10
D20995 N20995 0 diode
R20996 N20995 N20996 10
D20996 N20996 0 diode
R20997 N20996 N20997 10
D20997 N20997 0 diode
R20998 N20997 N20998 10
D20998 N20998 0 diode
R20999 N20998 N20999 10
D20999 N20999 0 diode
R21000 N20999 N21000 10
D21000 N21000 0 diode
R21001 N21000 N21001 10
D21001 N21001 0 diode
R21002 N21001 N21002 10
D21002 N21002 0 diode
R21003 N21002 N21003 10
D21003 N21003 0 diode
R21004 N21003 N21004 10
D21004 N21004 0 diode
R21005 N21004 N21005 10
D21005 N21005 0 diode
R21006 N21005 N21006 10
D21006 N21006 0 diode
R21007 N21006 N21007 10
D21007 N21007 0 diode
R21008 N21007 N21008 10
D21008 N21008 0 diode
R21009 N21008 N21009 10
D21009 N21009 0 diode
R21010 N21009 N21010 10
D21010 N21010 0 diode
R21011 N21010 N21011 10
D21011 N21011 0 diode
R21012 N21011 N21012 10
D21012 N21012 0 diode
R21013 N21012 N21013 10
D21013 N21013 0 diode
R21014 N21013 N21014 10
D21014 N21014 0 diode
R21015 N21014 N21015 10
D21015 N21015 0 diode
R21016 N21015 N21016 10
D21016 N21016 0 diode
R21017 N21016 N21017 10
D21017 N21017 0 diode
R21018 N21017 N21018 10
D21018 N21018 0 diode
R21019 N21018 N21019 10
D21019 N21019 0 diode
R21020 N21019 N21020 10
D21020 N21020 0 diode
R21021 N21020 N21021 10
D21021 N21021 0 diode
R21022 N21021 N21022 10
D21022 N21022 0 diode
R21023 N21022 N21023 10
D21023 N21023 0 diode
R21024 N21023 N21024 10
D21024 N21024 0 diode
R21025 N21024 N21025 10
D21025 N21025 0 diode
R21026 N21025 N21026 10
D21026 N21026 0 diode
R21027 N21026 N21027 10
D21027 N21027 0 diode
R21028 N21027 N21028 10
D21028 N21028 0 diode
R21029 N21028 N21029 10
D21029 N21029 0 diode
R21030 N21029 N21030 10
D21030 N21030 0 diode
R21031 N21030 N21031 10
D21031 N21031 0 diode
R21032 N21031 N21032 10
D21032 N21032 0 diode
R21033 N21032 N21033 10
D21033 N21033 0 diode
R21034 N21033 N21034 10
D21034 N21034 0 diode
R21035 N21034 N21035 10
D21035 N21035 0 diode
R21036 N21035 N21036 10
D21036 N21036 0 diode
R21037 N21036 N21037 10
D21037 N21037 0 diode
R21038 N21037 N21038 10
D21038 N21038 0 diode
R21039 N21038 N21039 10
D21039 N21039 0 diode
R21040 N21039 N21040 10
D21040 N21040 0 diode
R21041 N21040 N21041 10
D21041 N21041 0 diode
R21042 N21041 N21042 10
D21042 N21042 0 diode
R21043 N21042 N21043 10
D21043 N21043 0 diode
R21044 N21043 N21044 10
D21044 N21044 0 diode
R21045 N21044 N21045 10
D21045 N21045 0 diode
R21046 N21045 N21046 10
D21046 N21046 0 diode
R21047 N21046 N21047 10
D21047 N21047 0 diode
R21048 N21047 N21048 10
D21048 N21048 0 diode
R21049 N21048 N21049 10
D21049 N21049 0 diode
R21050 N21049 N21050 10
D21050 N21050 0 diode
R21051 N21050 N21051 10
D21051 N21051 0 diode
R21052 N21051 N21052 10
D21052 N21052 0 diode
R21053 N21052 N21053 10
D21053 N21053 0 diode
R21054 N21053 N21054 10
D21054 N21054 0 diode
R21055 N21054 N21055 10
D21055 N21055 0 diode
R21056 N21055 N21056 10
D21056 N21056 0 diode
R21057 N21056 N21057 10
D21057 N21057 0 diode
R21058 N21057 N21058 10
D21058 N21058 0 diode
R21059 N21058 N21059 10
D21059 N21059 0 diode
R21060 N21059 N21060 10
D21060 N21060 0 diode
R21061 N21060 N21061 10
D21061 N21061 0 diode
R21062 N21061 N21062 10
D21062 N21062 0 diode
R21063 N21062 N21063 10
D21063 N21063 0 diode
R21064 N21063 N21064 10
D21064 N21064 0 diode
R21065 N21064 N21065 10
D21065 N21065 0 diode
R21066 N21065 N21066 10
D21066 N21066 0 diode
R21067 N21066 N21067 10
D21067 N21067 0 diode
R21068 N21067 N21068 10
D21068 N21068 0 diode
R21069 N21068 N21069 10
D21069 N21069 0 diode
R21070 N21069 N21070 10
D21070 N21070 0 diode
R21071 N21070 N21071 10
D21071 N21071 0 diode
R21072 N21071 N21072 10
D21072 N21072 0 diode
R21073 N21072 N21073 10
D21073 N21073 0 diode
R21074 N21073 N21074 10
D21074 N21074 0 diode
R21075 N21074 N21075 10
D21075 N21075 0 diode
R21076 N21075 N21076 10
D21076 N21076 0 diode
R21077 N21076 N21077 10
D21077 N21077 0 diode
R21078 N21077 N21078 10
D21078 N21078 0 diode
R21079 N21078 N21079 10
D21079 N21079 0 diode
R21080 N21079 N21080 10
D21080 N21080 0 diode
R21081 N21080 N21081 10
D21081 N21081 0 diode
R21082 N21081 N21082 10
D21082 N21082 0 diode
R21083 N21082 N21083 10
D21083 N21083 0 diode
R21084 N21083 N21084 10
D21084 N21084 0 diode
R21085 N21084 N21085 10
D21085 N21085 0 diode
R21086 N21085 N21086 10
D21086 N21086 0 diode
R21087 N21086 N21087 10
D21087 N21087 0 diode
R21088 N21087 N21088 10
D21088 N21088 0 diode
R21089 N21088 N21089 10
D21089 N21089 0 diode
R21090 N21089 N21090 10
D21090 N21090 0 diode
R21091 N21090 N21091 10
D21091 N21091 0 diode
R21092 N21091 N21092 10
D21092 N21092 0 diode
R21093 N21092 N21093 10
D21093 N21093 0 diode
R21094 N21093 N21094 10
D21094 N21094 0 diode
R21095 N21094 N21095 10
D21095 N21095 0 diode
R21096 N21095 N21096 10
D21096 N21096 0 diode
R21097 N21096 N21097 10
D21097 N21097 0 diode
R21098 N21097 N21098 10
D21098 N21098 0 diode
R21099 N21098 N21099 10
D21099 N21099 0 diode
R21100 N21099 N21100 10
D21100 N21100 0 diode
R21101 N21100 N21101 10
D21101 N21101 0 diode
R21102 N21101 N21102 10
D21102 N21102 0 diode
R21103 N21102 N21103 10
D21103 N21103 0 diode
R21104 N21103 N21104 10
D21104 N21104 0 diode
R21105 N21104 N21105 10
D21105 N21105 0 diode
R21106 N21105 N21106 10
D21106 N21106 0 diode
R21107 N21106 N21107 10
D21107 N21107 0 diode
R21108 N21107 N21108 10
D21108 N21108 0 diode
R21109 N21108 N21109 10
D21109 N21109 0 diode
R21110 N21109 N21110 10
D21110 N21110 0 diode
R21111 N21110 N21111 10
D21111 N21111 0 diode
R21112 N21111 N21112 10
D21112 N21112 0 diode
R21113 N21112 N21113 10
D21113 N21113 0 diode
R21114 N21113 N21114 10
D21114 N21114 0 diode
R21115 N21114 N21115 10
D21115 N21115 0 diode
R21116 N21115 N21116 10
D21116 N21116 0 diode
R21117 N21116 N21117 10
D21117 N21117 0 diode
R21118 N21117 N21118 10
D21118 N21118 0 diode
R21119 N21118 N21119 10
D21119 N21119 0 diode
R21120 N21119 N21120 10
D21120 N21120 0 diode
R21121 N21120 N21121 10
D21121 N21121 0 diode
R21122 N21121 N21122 10
D21122 N21122 0 diode
R21123 N21122 N21123 10
D21123 N21123 0 diode
R21124 N21123 N21124 10
D21124 N21124 0 diode
R21125 N21124 N21125 10
D21125 N21125 0 diode
R21126 N21125 N21126 10
D21126 N21126 0 diode
R21127 N21126 N21127 10
D21127 N21127 0 diode
R21128 N21127 N21128 10
D21128 N21128 0 diode
R21129 N21128 N21129 10
D21129 N21129 0 diode
R21130 N21129 N21130 10
D21130 N21130 0 diode
R21131 N21130 N21131 10
D21131 N21131 0 diode
R21132 N21131 N21132 10
D21132 N21132 0 diode
R21133 N21132 N21133 10
D21133 N21133 0 diode
R21134 N21133 N21134 10
D21134 N21134 0 diode
R21135 N21134 N21135 10
D21135 N21135 0 diode
R21136 N21135 N21136 10
D21136 N21136 0 diode
R21137 N21136 N21137 10
D21137 N21137 0 diode
R21138 N21137 N21138 10
D21138 N21138 0 diode
R21139 N21138 N21139 10
D21139 N21139 0 diode
R21140 N21139 N21140 10
D21140 N21140 0 diode
R21141 N21140 N21141 10
D21141 N21141 0 diode
R21142 N21141 N21142 10
D21142 N21142 0 diode
R21143 N21142 N21143 10
D21143 N21143 0 diode
R21144 N21143 N21144 10
D21144 N21144 0 diode
R21145 N21144 N21145 10
D21145 N21145 0 diode
R21146 N21145 N21146 10
D21146 N21146 0 diode
R21147 N21146 N21147 10
D21147 N21147 0 diode
R21148 N21147 N21148 10
D21148 N21148 0 diode
R21149 N21148 N21149 10
D21149 N21149 0 diode
R21150 N21149 N21150 10
D21150 N21150 0 diode
R21151 N21150 N21151 10
D21151 N21151 0 diode
R21152 N21151 N21152 10
D21152 N21152 0 diode
R21153 N21152 N21153 10
D21153 N21153 0 diode
R21154 N21153 N21154 10
D21154 N21154 0 diode
R21155 N21154 N21155 10
D21155 N21155 0 diode
R21156 N21155 N21156 10
D21156 N21156 0 diode
R21157 N21156 N21157 10
D21157 N21157 0 diode
R21158 N21157 N21158 10
D21158 N21158 0 diode
R21159 N21158 N21159 10
D21159 N21159 0 diode
R21160 N21159 N21160 10
D21160 N21160 0 diode
R21161 N21160 N21161 10
D21161 N21161 0 diode
R21162 N21161 N21162 10
D21162 N21162 0 diode
R21163 N21162 N21163 10
D21163 N21163 0 diode
R21164 N21163 N21164 10
D21164 N21164 0 diode
R21165 N21164 N21165 10
D21165 N21165 0 diode
R21166 N21165 N21166 10
D21166 N21166 0 diode
R21167 N21166 N21167 10
D21167 N21167 0 diode
R21168 N21167 N21168 10
D21168 N21168 0 diode
R21169 N21168 N21169 10
D21169 N21169 0 diode
R21170 N21169 N21170 10
D21170 N21170 0 diode
R21171 N21170 N21171 10
D21171 N21171 0 diode
R21172 N21171 N21172 10
D21172 N21172 0 diode
R21173 N21172 N21173 10
D21173 N21173 0 diode
R21174 N21173 N21174 10
D21174 N21174 0 diode
R21175 N21174 N21175 10
D21175 N21175 0 diode
R21176 N21175 N21176 10
D21176 N21176 0 diode
R21177 N21176 N21177 10
D21177 N21177 0 diode
R21178 N21177 N21178 10
D21178 N21178 0 diode
R21179 N21178 N21179 10
D21179 N21179 0 diode
R21180 N21179 N21180 10
D21180 N21180 0 diode
R21181 N21180 N21181 10
D21181 N21181 0 diode
R21182 N21181 N21182 10
D21182 N21182 0 diode
R21183 N21182 N21183 10
D21183 N21183 0 diode
R21184 N21183 N21184 10
D21184 N21184 0 diode
R21185 N21184 N21185 10
D21185 N21185 0 diode
R21186 N21185 N21186 10
D21186 N21186 0 diode
R21187 N21186 N21187 10
D21187 N21187 0 diode
R21188 N21187 N21188 10
D21188 N21188 0 diode
R21189 N21188 N21189 10
D21189 N21189 0 diode
R21190 N21189 N21190 10
D21190 N21190 0 diode
R21191 N21190 N21191 10
D21191 N21191 0 diode
R21192 N21191 N21192 10
D21192 N21192 0 diode
R21193 N21192 N21193 10
D21193 N21193 0 diode
R21194 N21193 N21194 10
D21194 N21194 0 diode
R21195 N21194 N21195 10
D21195 N21195 0 diode
R21196 N21195 N21196 10
D21196 N21196 0 diode
R21197 N21196 N21197 10
D21197 N21197 0 diode
R21198 N21197 N21198 10
D21198 N21198 0 diode
R21199 N21198 N21199 10
D21199 N21199 0 diode
R21200 N21199 N21200 10
D21200 N21200 0 diode
R21201 N21200 N21201 10
D21201 N21201 0 diode
R21202 N21201 N21202 10
D21202 N21202 0 diode
R21203 N21202 N21203 10
D21203 N21203 0 diode
R21204 N21203 N21204 10
D21204 N21204 0 diode
R21205 N21204 N21205 10
D21205 N21205 0 diode
R21206 N21205 N21206 10
D21206 N21206 0 diode
R21207 N21206 N21207 10
D21207 N21207 0 diode
R21208 N21207 N21208 10
D21208 N21208 0 diode
R21209 N21208 N21209 10
D21209 N21209 0 diode
R21210 N21209 N21210 10
D21210 N21210 0 diode
R21211 N21210 N21211 10
D21211 N21211 0 diode
R21212 N21211 N21212 10
D21212 N21212 0 diode
R21213 N21212 N21213 10
D21213 N21213 0 diode
R21214 N21213 N21214 10
D21214 N21214 0 diode
R21215 N21214 N21215 10
D21215 N21215 0 diode
R21216 N21215 N21216 10
D21216 N21216 0 diode
R21217 N21216 N21217 10
D21217 N21217 0 diode
R21218 N21217 N21218 10
D21218 N21218 0 diode
R21219 N21218 N21219 10
D21219 N21219 0 diode
R21220 N21219 N21220 10
D21220 N21220 0 diode
R21221 N21220 N21221 10
D21221 N21221 0 diode
R21222 N21221 N21222 10
D21222 N21222 0 diode
R21223 N21222 N21223 10
D21223 N21223 0 diode
R21224 N21223 N21224 10
D21224 N21224 0 diode
R21225 N21224 N21225 10
D21225 N21225 0 diode
R21226 N21225 N21226 10
D21226 N21226 0 diode
R21227 N21226 N21227 10
D21227 N21227 0 diode
R21228 N21227 N21228 10
D21228 N21228 0 diode
R21229 N21228 N21229 10
D21229 N21229 0 diode
R21230 N21229 N21230 10
D21230 N21230 0 diode
R21231 N21230 N21231 10
D21231 N21231 0 diode
R21232 N21231 N21232 10
D21232 N21232 0 diode
R21233 N21232 N21233 10
D21233 N21233 0 diode
R21234 N21233 N21234 10
D21234 N21234 0 diode
R21235 N21234 N21235 10
D21235 N21235 0 diode
R21236 N21235 N21236 10
D21236 N21236 0 diode
R21237 N21236 N21237 10
D21237 N21237 0 diode
R21238 N21237 N21238 10
D21238 N21238 0 diode
R21239 N21238 N21239 10
D21239 N21239 0 diode
R21240 N21239 N21240 10
D21240 N21240 0 diode
R21241 N21240 N21241 10
D21241 N21241 0 diode
R21242 N21241 N21242 10
D21242 N21242 0 diode
R21243 N21242 N21243 10
D21243 N21243 0 diode
R21244 N21243 N21244 10
D21244 N21244 0 diode
R21245 N21244 N21245 10
D21245 N21245 0 diode
R21246 N21245 N21246 10
D21246 N21246 0 diode
R21247 N21246 N21247 10
D21247 N21247 0 diode
R21248 N21247 N21248 10
D21248 N21248 0 diode
R21249 N21248 N21249 10
D21249 N21249 0 diode
R21250 N21249 N21250 10
D21250 N21250 0 diode
R21251 N21250 N21251 10
D21251 N21251 0 diode
R21252 N21251 N21252 10
D21252 N21252 0 diode
R21253 N21252 N21253 10
D21253 N21253 0 diode
R21254 N21253 N21254 10
D21254 N21254 0 diode
R21255 N21254 N21255 10
D21255 N21255 0 diode
R21256 N21255 N21256 10
D21256 N21256 0 diode
R21257 N21256 N21257 10
D21257 N21257 0 diode
R21258 N21257 N21258 10
D21258 N21258 0 diode
R21259 N21258 N21259 10
D21259 N21259 0 diode
R21260 N21259 N21260 10
D21260 N21260 0 diode
R21261 N21260 N21261 10
D21261 N21261 0 diode
R21262 N21261 N21262 10
D21262 N21262 0 diode
R21263 N21262 N21263 10
D21263 N21263 0 diode
R21264 N21263 N21264 10
D21264 N21264 0 diode
R21265 N21264 N21265 10
D21265 N21265 0 diode
R21266 N21265 N21266 10
D21266 N21266 0 diode
R21267 N21266 N21267 10
D21267 N21267 0 diode
R21268 N21267 N21268 10
D21268 N21268 0 diode
R21269 N21268 N21269 10
D21269 N21269 0 diode
R21270 N21269 N21270 10
D21270 N21270 0 diode
R21271 N21270 N21271 10
D21271 N21271 0 diode
R21272 N21271 N21272 10
D21272 N21272 0 diode
R21273 N21272 N21273 10
D21273 N21273 0 diode
R21274 N21273 N21274 10
D21274 N21274 0 diode
R21275 N21274 N21275 10
D21275 N21275 0 diode
R21276 N21275 N21276 10
D21276 N21276 0 diode
R21277 N21276 N21277 10
D21277 N21277 0 diode
R21278 N21277 N21278 10
D21278 N21278 0 diode
R21279 N21278 N21279 10
D21279 N21279 0 diode
R21280 N21279 N21280 10
D21280 N21280 0 diode
R21281 N21280 N21281 10
D21281 N21281 0 diode
R21282 N21281 N21282 10
D21282 N21282 0 diode
R21283 N21282 N21283 10
D21283 N21283 0 diode
R21284 N21283 N21284 10
D21284 N21284 0 diode
R21285 N21284 N21285 10
D21285 N21285 0 diode
R21286 N21285 N21286 10
D21286 N21286 0 diode
R21287 N21286 N21287 10
D21287 N21287 0 diode
R21288 N21287 N21288 10
D21288 N21288 0 diode
R21289 N21288 N21289 10
D21289 N21289 0 diode
R21290 N21289 N21290 10
D21290 N21290 0 diode
R21291 N21290 N21291 10
D21291 N21291 0 diode
R21292 N21291 N21292 10
D21292 N21292 0 diode
R21293 N21292 N21293 10
D21293 N21293 0 diode
R21294 N21293 N21294 10
D21294 N21294 0 diode
R21295 N21294 N21295 10
D21295 N21295 0 diode
R21296 N21295 N21296 10
D21296 N21296 0 diode
R21297 N21296 N21297 10
D21297 N21297 0 diode
R21298 N21297 N21298 10
D21298 N21298 0 diode
R21299 N21298 N21299 10
D21299 N21299 0 diode
R21300 N21299 N21300 10
D21300 N21300 0 diode
R21301 N21300 N21301 10
D21301 N21301 0 diode
R21302 N21301 N21302 10
D21302 N21302 0 diode
R21303 N21302 N21303 10
D21303 N21303 0 diode
R21304 N21303 N21304 10
D21304 N21304 0 diode
R21305 N21304 N21305 10
D21305 N21305 0 diode
R21306 N21305 N21306 10
D21306 N21306 0 diode
R21307 N21306 N21307 10
D21307 N21307 0 diode
R21308 N21307 N21308 10
D21308 N21308 0 diode
R21309 N21308 N21309 10
D21309 N21309 0 diode
R21310 N21309 N21310 10
D21310 N21310 0 diode
R21311 N21310 N21311 10
D21311 N21311 0 diode
R21312 N21311 N21312 10
D21312 N21312 0 diode
R21313 N21312 N21313 10
D21313 N21313 0 diode
R21314 N21313 N21314 10
D21314 N21314 0 diode
R21315 N21314 N21315 10
D21315 N21315 0 diode
R21316 N21315 N21316 10
D21316 N21316 0 diode
R21317 N21316 N21317 10
D21317 N21317 0 diode
R21318 N21317 N21318 10
D21318 N21318 0 diode
R21319 N21318 N21319 10
D21319 N21319 0 diode
R21320 N21319 N21320 10
D21320 N21320 0 diode
R21321 N21320 N21321 10
D21321 N21321 0 diode
R21322 N21321 N21322 10
D21322 N21322 0 diode
R21323 N21322 N21323 10
D21323 N21323 0 diode
R21324 N21323 N21324 10
D21324 N21324 0 diode
R21325 N21324 N21325 10
D21325 N21325 0 diode
R21326 N21325 N21326 10
D21326 N21326 0 diode
R21327 N21326 N21327 10
D21327 N21327 0 diode
R21328 N21327 N21328 10
D21328 N21328 0 diode
R21329 N21328 N21329 10
D21329 N21329 0 diode
R21330 N21329 N21330 10
D21330 N21330 0 diode
R21331 N21330 N21331 10
D21331 N21331 0 diode
R21332 N21331 N21332 10
D21332 N21332 0 diode
R21333 N21332 N21333 10
D21333 N21333 0 diode
R21334 N21333 N21334 10
D21334 N21334 0 diode
R21335 N21334 N21335 10
D21335 N21335 0 diode
R21336 N21335 N21336 10
D21336 N21336 0 diode
R21337 N21336 N21337 10
D21337 N21337 0 diode
R21338 N21337 N21338 10
D21338 N21338 0 diode
R21339 N21338 N21339 10
D21339 N21339 0 diode
R21340 N21339 N21340 10
D21340 N21340 0 diode
R21341 N21340 N21341 10
D21341 N21341 0 diode
R21342 N21341 N21342 10
D21342 N21342 0 diode
R21343 N21342 N21343 10
D21343 N21343 0 diode
R21344 N21343 N21344 10
D21344 N21344 0 diode
R21345 N21344 N21345 10
D21345 N21345 0 diode
R21346 N21345 N21346 10
D21346 N21346 0 diode
R21347 N21346 N21347 10
D21347 N21347 0 diode
R21348 N21347 N21348 10
D21348 N21348 0 diode
R21349 N21348 N21349 10
D21349 N21349 0 diode
R21350 N21349 N21350 10
D21350 N21350 0 diode
R21351 N21350 N21351 10
D21351 N21351 0 diode
R21352 N21351 N21352 10
D21352 N21352 0 diode
R21353 N21352 N21353 10
D21353 N21353 0 diode
R21354 N21353 N21354 10
D21354 N21354 0 diode
R21355 N21354 N21355 10
D21355 N21355 0 diode
R21356 N21355 N21356 10
D21356 N21356 0 diode
R21357 N21356 N21357 10
D21357 N21357 0 diode
R21358 N21357 N21358 10
D21358 N21358 0 diode
R21359 N21358 N21359 10
D21359 N21359 0 diode
R21360 N21359 N21360 10
D21360 N21360 0 diode
R21361 N21360 N21361 10
D21361 N21361 0 diode
R21362 N21361 N21362 10
D21362 N21362 0 diode
R21363 N21362 N21363 10
D21363 N21363 0 diode
R21364 N21363 N21364 10
D21364 N21364 0 diode
R21365 N21364 N21365 10
D21365 N21365 0 diode
R21366 N21365 N21366 10
D21366 N21366 0 diode
R21367 N21366 N21367 10
D21367 N21367 0 diode
R21368 N21367 N21368 10
D21368 N21368 0 diode
R21369 N21368 N21369 10
D21369 N21369 0 diode
R21370 N21369 N21370 10
D21370 N21370 0 diode
R21371 N21370 N21371 10
D21371 N21371 0 diode
R21372 N21371 N21372 10
D21372 N21372 0 diode
R21373 N21372 N21373 10
D21373 N21373 0 diode
R21374 N21373 N21374 10
D21374 N21374 0 diode
R21375 N21374 N21375 10
D21375 N21375 0 diode
R21376 N21375 N21376 10
D21376 N21376 0 diode
R21377 N21376 N21377 10
D21377 N21377 0 diode
R21378 N21377 N21378 10
D21378 N21378 0 diode
R21379 N21378 N21379 10
D21379 N21379 0 diode
R21380 N21379 N21380 10
D21380 N21380 0 diode
R21381 N21380 N21381 10
D21381 N21381 0 diode
R21382 N21381 N21382 10
D21382 N21382 0 diode
R21383 N21382 N21383 10
D21383 N21383 0 diode
R21384 N21383 N21384 10
D21384 N21384 0 diode
R21385 N21384 N21385 10
D21385 N21385 0 diode
R21386 N21385 N21386 10
D21386 N21386 0 diode
R21387 N21386 N21387 10
D21387 N21387 0 diode
R21388 N21387 N21388 10
D21388 N21388 0 diode
R21389 N21388 N21389 10
D21389 N21389 0 diode
R21390 N21389 N21390 10
D21390 N21390 0 diode
R21391 N21390 N21391 10
D21391 N21391 0 diode
R21392 N21391 N21392 10
D21392 N21392 0 diode
R21393 N21392 N21393 10
D21393 N21393 0 diode
R21394 N21393 N21394 10
D21394 N21394 0 diode
R21395 N21394 N21395 10
D21395 N21395 0 diode
R21396 N21395 N21396 10
D21396 N21396 0 diode
R21397 N21396 N21397 10
D21397 N21397 0 diode
R21398 N21397 N21398 10
D21398 N21398 0 diode
R21399 N21398 N21399 10
D21399 N21399 0 diode
R21400 N21399 N21400 10
D21400 N21400 0 diode
R21401 N21400 N21401 10
D21401 N21401 0 diode
R21402 N21401 N21402 10
D21402 N21402 0 diode
R21403 N21402 N21403 10
D21403 N21403 0 diode
R21404 N21403 N21404 10
D21404 N21404 0 diode
R21405 N21404 N21405 10
D21405 N21405 0 diode
R21406 N21405 N21406 10
D21406 N21406 0 diode
R21407 N21406 N21407 10
D21407 N21407 0 diode
R21408 N21407 N21408 10
D21408 N21408 0 diode
R21409 N21408 N21409 10
D21409 N21409 0 diode
R21410 N21409 N21410 10
D21410 N21410 0 diode
R21411 N21410 N21411 10
D21411 N21411 0 diode
R21412 N21411 N21412 10
D21412 N21412 0 diode
R21413 N21412 N21413 10
D21413 N21413 0 diode
R21414 N21413 N21414 10
D21414 N21414 0 diode
R21415 N21414 N21415 10
D21415 N21415 0 diode
R21416 N21415 N21416 10
D21416 N21416 0 diode
R21417 N21416 N21417 10
D21417 N21417 0 diode
R21418 N21417 N21418 10
D21418 N21418 0 diode
R21419 N21418 N21419 10
D21419 N21419 0 diode
R21420 N21419 N21420 10
D21420 N21420 0 diode
R21421 N21420 N21421 10
D21421 N21421 0 diode
R21422 N21421 N21422 10
D21422 N21422 0 diode
R21423 N21422 N21423 10
D21423 N21423 0 diode
R21424 N21423 N21424 10
D21424 N21424 0 diode
R21425 N21424 N21425 10
D21425 N21425 0 diode
R21426 N21425 N21426 10
D21426 N21426 0 diode
R21427 N21426 N21427 10
D21427 N21427 0 diode
R21428 N21427 N21428 10
D21428 N21428 0 diode
R21429 N21428 N21429 10
D21429 N21429 0 diode
R21430 N21429 N21430 10
D21430 N21430 0 diode
R21431 N21430 N21431 10
D21431 N21431 0 diode
R21432 N21431 N21432 10
D21432 N21432 0 diode
R21433 N21432 N21433 10
D21433 N21433 0 diode
R21434 N21433 N21434 10
D21434 N21434 0 diode
R21435 N21434 N21435 10
D21435 N21435 0 diode
R21436 N21435 N21436 10
D21436 N21436 0 diode
R21437 N21436 N21437 10
D21437 N21437 0 diode
R21438 N21437 N21438 10
D21438 N21438 0 diode
R21439 N21438 N21439 10
D21439 N21439 0 diode
R21440 N21439 N21440 10
D21440 N21440 0 diode
R21441 N21440 N21441 10
D21441 N21441 0 diode
R21442 N21441 N21442 10
D21442 N21442 0 diode
R21443 N21442 N21443 10
D21443 N21443 0 diode
R21444 N21443 N21444 10
D21444 N21444 0 diode
R21445 N21444 N21445 10
D21445 N21445 0 diode
R21446 N21445 N21446 10
D21446 N21446 0 diode
R21447 N21446 N21447 10
D21447 N21447 0 diode
R21448 N21447 N21448 10
D21448 N21448 0 diode
R21449 N21448 N21449 10
D21449 N21449 0 diode
R21450 N21449 N21450 10
D21450 N21450 0 diode
R21451 N21450 N21451 10
D21451 N21451 0 diode
R21452 N21451 N21452 10
D21452 N21452 0 diode
R21453 N21452 N21453 10
D21453 N21453 0 diode
R21454 N21453 N21454 10
D21454 N21454 0 diode
R21455 N21454 N21455 10
D21455 N21455 0 diode
R21456 N21455 N21456 10
D21456 N21456 0 diode
R21457 N21456 N21457 10
D21457 N21457 0 diode
R21458 N21457 N21458 10
D21458 N21458 0 diode
R21459 N21458 N21459 10
D21459 N21459 0 diode
R21460 N21459 N21460 10
D21460 N21460 0 diode
R21461 N21460 N21461 10
D21461 N21461 0 diode
R21462 N21461 N21462 10
D21462 N21462 0 diode
R21463 N21462 N21463 10
D21463 N21463 0 diode
R21464 N21463 N21464 10
D21464 N21464 0 diode
R21465 N21464 N21465 10
D21465 N21465 0 diode
R21466 N21465 N21466 10
D21466 N21466 0 diode
R21467 N21466 N21467 10
D21467 N21467 0 diode
R21468 N21467 N21468 10
D21468 N21468 0 diode
R21469 N21468 N21469 10
D21469 N21469 0 diode
R21470 N21469 N21470 10
D21470 N21470 0 diode
R21471 N21470 N21471 10
D21471 N21471 0 diode
R21472 N21471 N21472 10
D21472 N21472 0 diode
R21473 N21472 N21473 10
D21473 N21473 0 diode
R21474 N21473 N21474 10
D21474 N21474 0 diode
R21475 N21474 N21475 10
D21475 N21475 0 diode
R21476 N21475 N21476 10
D21476 N21476 0 diode
R21477 N21476 N21477 10
D21477 N21477 0 diode
R21478 N21477 N21478 10
D21478 N21478 0 diode
R21479 N21478 N21479 10
D21479 N21479 0 diode
R21480 N21479 N21480 10
D21480 N21480 0 diode
R21481 N21480 N21481 10
D21481 N21481 0 diode
R21482 N21481 N21482 10
D21482 N21482 0 diode
R21483 N21482 N21483 10
D21483 N21483 0 diode
R21484 N21483 N21484 10
D21484 N21484 0 diode
R21485 N21484 N21485 10
D21485 N21485 0 diode
R21486 N21485 N21486 10
D21486 N21486 0 diode
R21487 N21486 N21487 10
D21487 N21487 0 diode
R21488 N21487 N21488 10
D21488 N21488 0 diode
R21489 N21488 N21489 10
D21489 N21489 0 diode
R21490 N21489 N21490 10
D21490 N21490 0 diode
R21491 N21490 N21491 10
D21491 N21491 0 diode
R21492 N21491 N21492 10
D21492 N21492 0 diode
R21493 N21492 N21493 10
D21493 N21493 0 diode
R21494 N21493 N21494 10
D21494 N21494 0 diode
R21495 N21494 N21495 10
D21495 N21495 0 diode
R21496 N21495 N21496 10
D21496 N21496 0 diode
R21497 N21496 N21497 10
D21497 N21497 0 diode
R21498 N21497 N21498 10
D21498 N21498 0 diode
R21499 N21498 N21499 10
D21499 N21499 0 diode
R21500 N21499 N21500 10
D21500 N21500 0 diode
R21501 N21500 N21501 10
D21501 N21501 0 diode
R21502 N21501 N21502 10
D21502 N21502 0 diode
R21503 N21502 N21503 10
D21503 N21503 0 diode
R21504 N21503 N21504 10
D21504 N21504 0 diode
R21505 N21504 N21505 10
D21505 N21505 0 diode
R21506 N21505 N21506 10
D21506 N21506 0 diode
R21507 N21506 N21507 10
D21507 N21507 0 diode
R21508 N21507 N21508 10
D21508 N21508 0 diode
R21509 N21508 N21509 10
D21509 N21509 0 diode
R21510 N21509 N21510 10
D21510 N21510 0 diode
R21511 N21510 N21511 10
D21511 N21511 0 diode
R21512 N21511 N21512 10
D21512 N21512 0 diode
R21513 N21512 N21513 10
D21513 N21513 0 diode
R21514 N21513 N21514 10
D21514 N21514 0 diode
R21515 N21514 N21515 10
D21515 N21515 0 diode
R21516 N21515 N21516 10
D21516 N21516 0 diode
R21517 N21516 N21517 10
D21517 N21517 0 diode
R21518 N21517 N21518 10
D21518 N21518 0 diode
R21519 N21518 N21519 10
D21519 N21519 0 diode
R21520 N21519 N21520 10
D21520 N21520 0 diode
R21521 N21520 N21521 10
D21521 N21521 0 diode
R21522 N21521 N21522 10
D21522 N21522 0 diode
R21523 N21522 N21523 10
D21523 N21523 0 diode
R21524 N21523 N21524 10
D21524 N21524 0 diode
R21525 N21524 N21525 10
D21525 N21525 0 diode
R21526 N21525 N21526 10
D21526 N21526 0 diode
R21527 N21526 N21527 10
D21527 N21527 0 diode
R21528 N21527 N21528 10
D21528 N21528 0 diode
R21529 N21528 N21529 10
D21529 N21529 0 diode
R21530 N21529 N21530 10
D21530 N21530 0 diode
R21531 N21530 N21531 10
D21531 N21531 0 diode
R21532 N21531 N21532 10
D21532 N21532 0 diode
R21533 N21532 N21533 10
D21533 N21533 0 diode
R21534 N21533 N21534 10
D21534 N21534 0 diode
R21535 N21534 N21535 10
D21535 N21535 0 diode
R21536 N21535 N21536 10
D21536 N21536 0 diode
R21537 N21536 N21537 10
D21537 N21537 0 diode
R21538 N21537 N21538 10
D21538 N21538 0 diode
R21539 N21538 N21539 10
D21539 N21539 0 diode
R21540 N21539 N21540 10
D21540 N21540 0 diode
R21541 N21540 N21541 10
D21541 N21541 0 diode
R21542 N21541 N21542 10
D21542 N21542 0 diode
R21543 N21542 N21543 10
D21543 N21543 0 diode
R21544 N21543 N21544 10
D21544 N21544 0 diode
R21545 N21544 N21545 10
D21545 N21545 0 diode
R21546 N21545 N21546 10
D21546 N21546 0 diode
R21547 N21546 N21547 10
D21547 N21547 0 diode
R21548 N21547 N21548 10
D21548 N21548 0 diode
R21549 N21548 N21549 10
D21549 N21549 0 diode
R21550 N21549 N21550 10
D21550 N21550 0 diode
R21551 N21550 N21551 10
D21551 N21551 0 diode
R21552 N21551 N21552 10
D21552 N21552 0 diode
R21553 N21552 N21553 10
D21553 N21553 0 diode
R21554 N21553 N21554 10
D21554 N21554 0 diode
R21555 N21554 N21555 10
D21555 N21555 0 diode
R21556 N21555 N21556 10
D21556 N21556 0 diode
R21557 N21556 N21557 10
D21557 N21557 0 diode
R21558 N21557 N21558 10
D21558 N21558 0 diode
R21559 N21558 N21559 10
D21559 N21559 0 diode
R21560 N21559 N21560 10
D21560 N21560 0 diode
R21561 N21560 N21561 10
D21561 N21561 0 diode
R21562 N21561 N21562 10
D21562 N21562 0 diode
R21563 N21562 N21563 10
D21563 N21563 0 diode
R21564 N21563 N21564 10
D21564 N21564 0 diode
R21565 N21564 N21565 10
D21565 N21565 0 diode
R21566 N21565 N21566 10
D21566 N21566 0 diode
R21567 N21566 N21567 10
D21567 N21567 0 diode
R21568 N21567 N21568 10
D21568 N21568 0 diode
R21569 N21568 N21569 10
D21569 N21569 0 diode
R21570 N21569 N21570 10
D21570 N21570 0 diode
R21571 N21570 N21571 10
D21571 N21571 0 diode
R21572 N21571 N21572 10
D21572 N21572 0 diode
R21573 N21572 N21573 10
D21573 N21573 0 diode
R21574 N21573 N21574 10
D21574 N21574 0 diode
R21575 N21574 N21575 10
D21575 N21575 0 diode
R21576 N21575 N21576 10
D21576 N21576 0 diode
R21577 N21576 N21577 10
D21577 N21577 0 diode
R21578 N21577 N21578 10
D21578 N21578 0 diode
R21579 N21578 N21579 10
D21579 N21579 0 diode
R21580 N21579 N21580 10
D21580 N21580 0 diode
R21581 N21580 N21581 10
D21581 N21581 0 diode
R21582 N21581 N21582 10
D21582 N21582 0 diode
R21583 N21582 N21583 10
D21583 N21583 0 diode
R21584 N21583 N21584 10
D21584 N21584 0 diode
R21585 N21584 N21585 10
D21585 N21585 0 diode
R21586 N21585 N21586 10
D21586 N21586 0 diode
R21587 N21586 N21587 10
D21587 N21587 0 diode
R21588 N21587 N21588 10
D21588 N21588 0 diode
R21589 N21588 N21589 10
D21589 N21589 0 diode
R21590 N21589 N21590 10
D21590 N21590 0 diode
R21591 N21590 N21591 10
D21591 N21591 0 diode
R21592 N21591 N21592 10
D21592 N21592 0 diode
R21593 N21592 N21593 10
D21593 N21593 0 diode
R21594 N21593 N21594 10
D21594 N21594 0 diode
R21595 N21594 N21595 10
D21595 N21595 0 diode
R21596 N21595 N21596 10
D21596 N21596 0 diode
R21597 N21596 N21597 10
D21597 N21597 0 diode
R21598 N21597 N21598 10
D21598 N21598 0 diode
R21599 N21598 N21599 10
D21599 N21599 0 diode
R21600 N21599 N21600 10
D21600 N21600 0 diode
R21601 N21600 N21601 10
D21601 N21601 0 diode
R21602 N21601 N21602 10
D21602 N21602 0 diode
R21603 N21602 N21603 10
D21603 N21603 0 diode
R21604 N21603 N21604 10
D21604 N21604 0 diode
R21605 N21604 N21605 10
D21605 N21605 0 diode
R21606 N21605 N21606 10
D21606 N21606 0 diode
R21607 N21606 N21607 10
D21607 N21607 0 diode
R21608 N21607 N21608 10
D21608 N21608 0 diode
R21609 N21608 N21609 10
D21609 N21609 0 diode
R21610 N21609 N21610 10
D21610 N21610 0 diode
R21611 N21610 N21611 10
D21611 N21611 0 diode
R21612 N21611 N21612 10
D21612 N21612 0 diode
R21613 N21612 N21613 10
D21613 N21613 0 diode
R21614 N21613 N21614 10
D21614 N21614 0 diode
R21615 N21614 N21615 10
D21615 N21615 0 diode
R21616 N21615 N21616 10
D21616 N21616 0 diode
R21617 N21616 N21617 10
D21617 N21617 0 diode
R21618 N21617 N21618 10
D21618 N21618 0 diode
R21619 N21618 N21619 10
D21619 N21619 0 diode
R21620 N21619 N21620 10
D21620 N21620 0 diode
R21621 N21620 N21621 10
D21621 N21621 0 diode
R21622 N21621 N21622 10
D21622 N21622 0 diode
R21623 N21622 N21623 10
D21623 N21623 0 diode
R21624 N21623 N21624 10
D21624 N21624 0 diode
R21625 N21624 N21625 10
D21625 N21625 0 diode
R21626 N21625 N21626 10
D21626 N21626 0 diode
R21627 N21626 N21627 10
D21627 N21627 0 diode
R21628 N21627 N21628 10
D21628 N21628 0 diode
R21629 N21628 N21629 10
D21629 N21629 0 diode
R21630 N21629 N21630 10
D21630 N21630 0 diode
R21631 N21630 N21631 10
D21631 N21631 0 diode
R21632 N21631 N21632 10
D21632 N21632 0 diode
R21633 N21632 N21633 10
D21633 N21633 0 diode
R21634 N21633 N21634 10
D21634 N21634 0 diode
R21635 N21634 N21635 10
D21635 N21635 0 diode
R21636 N21635 N21636 10
D21636 N21636 0 diode
R21637 N21636 N21637 10
D21637 N21637 0 diode
R21638 N21637 N21638 10
D21638 N21638 0 diode
R21639 N21638 N21639 10
D21639 N21639 0 diode
R21640 N21639 N21640 10
D21640 N21640 0 diode
R21641 N21640 N21641 10
D21641 N21641 0 diode
R21642 N21641 N21642 10
D21642 N21642 0 diode
R21643 N21642 N21643 10
D21643 N21643 0 diode
R21644 N21643 N21644 10
D21644 N21644 0 diode
R21645 N21644 N21645 10
D21645 N21645 0 diode
R21646 N21645 N21646 10
D21646 N21646 0 diode
R21647 N21646 N21647 10
D21647 N21647 0 diode
R21648 N21647 N21648 10
D21648 N21648 0 diode
R21649 N21648 N21649 10
D21649 N21649 0 diode
R21650 N21649 N21650 10
D21650 N21650 0 diode
R21651 N21650 N21651 10
D21651 N21651 0 diode
R21652 N21651 N21652 10
D21652 N21652 0 diode
R21653 N21652 N21653 10
D21653 N21653 0 diode
R21654 N21653 N21654 10
D21654 N21654 0 diode
R21655 N21654 N21655 10
D21655 N21655 0 diode
R21656 N21655 N21656 10
D21656 N21656 0 diode
R21657 N21656 N21657 10
D21657 N21657 0 diode
R21658 N21657 N21658 10
D21658 N21658 0 diode
R21659 N21658 N21659 10
D21659 N21659 0 diode
R21660 N21659 N21660 10
D21660 N21660 0 diode
R21661 N21660 N21661 10
D21661 N21661 0 diode
R21662 N21661 N21662 10
D21662 N21662 0 diode
R21663 N21662 N21663 10
D21663 N21663 0 diode
R21664 N21663 N21664 10
D21664 N21664 0 diode
R21665 N21664 N21665 10
D21665 N21665 0 diode
R21666 N21665 N21666 10
D21666 N21666 0 diode
R21667 N21666 N21667 10
D21667 N21667 0 diode
R21668 N21667 N21668 10
D21668 N21668 0 diode
R21669 N21668 N21669 10
D21669 N21669 0 diode
R21670 N21669 N21670 10
D21670 N21670 0 diode
R21671 N21670 N21671 10
D21671 N21671 0 diode
R21672 N21671 N21672 10
D21672 N21672 0 diode
R21673 N21672 N21673 10
D21673 N21673 0 diode
R21674 N21673 N21674 10
D21674 N21674 0 diode
R21675 N21674 N21675 10
D21675 N21675 0 diode
R21676 N21675 N21676 10
D21676 N21676 0 diode
R21677 N21676 N21677 10
D21677 N21677 0 diode
R21678 N21677 N21678 10
D21678 N21678 0 diode
R21679 N21678 N21679 10
D21679 N21679 0 diode
R21680 N21679 N21680 10
D21680 N21680 0 diode
R21681 N21680 N21681 10
D21681 N21681 0 diode
R21682 N21681 N21682 10
D21682 N21682 0 diode
R21683 N21682 N21683 10
D21683 N21683 0 diode
R21684 N21683 N21684 10
D21684 N21684 0 diode
R21685 N21684 N21685 10
D21685 N21685 0 diode
R21686 N21685 N21686 10
D21686 N21686 0 diode
R21687 N21686 N21687 10
D21687 N21687 0 diode
R21688 N21687 N21688 10
D21688 N21688 0 diode
R21689 N21688 N21689 10
D21689 N21689 0 diode
R21690 N21689 N21690 10
D21690 N21690 0 diode
R21691 N21690 N21691 10
D21691 N21691 0 diode
R21692 N21691 N21692 10
D21692 N21692 0 diode
R21693 N21692 N21693 10
D21693 N21693 0 diode
R21694 N21693 N21694 10
D21694 N21694 0 diode
R21695 N21694 N21695 10
D21695 N21695 0 diode
R21696 N21695 N21696 10
D21696 N21696 0 diode
R21697 N21696 N21697 10
D21697 N21697 0 diode
R21698 N21697 N21698 10
D21698 N21698 0 diode
R21699 N21698 N21699 10
D21699 N21699 0 diode
R21700 N21699 N21700 10
D21700 N21700 0 diode
R21701 N21700 N21701 10
D21701 N21701 0 diode
R21702 N21701 N21702 10
D21702 N21702 0 diode
R21703 N21702 N21703 10
D21703 N21703 0 diode
R21704 N21703 N21704 10
D21704 N21704 0 diode
R21705 N21704 N21705 10
D21705 N21705 0 diode
R21706 N21705 N21706 10
D21706 N21706 0 diode
R21707 N21706 N21707 10
D21707 N21707 0 diode
R21708 N21707 N21708 10
D21708 N21708 0 diode
R21709 N21708 N21709 10
D21709 N21709 0 diode
R21710 N21709 N21710 10
D21710 N21710 0 diode
R21711 N21710 N21711 10
D21711 N21711 0 diode
R21712 N21711 N21712 10
D21712 N21712 0 diode
R21713 N21712 N21713 10
D21713 N21713 0 diode
R21714 N21713 N21714 10
D21714 N21714 0 diode
R21715 N21714 N21715 10
D21715 N21715 0 diode
R21716 N21715 N21716 10
D21716 N21716 0 diode
R21717 N21716 N21717 10
D21717 N21717 0 diode
R21718 N21717 N21718 10
D21718 N21718 0 diode
R21719 N21718 N21719 10
D21719 N21719 0 diode
R21720 N21719 N21720 10
D21720 N21720 0 diode
R21721 N21720 N21721 10
D21721 N21721 0 diode
R21722 N21721 N21722 10
D21722 N21722 0 diode
R21723 N21722 N21723 10
D21723 N21723 0 diode
R21724 N21723 N21724 10
D21724 N21724 0 diode
R21725 N21724 N21725 10
D21725 N21725 0 diode
R21726 N21725 N21726 10
D21726 N21726 0 diode
R21727 N21726 N21727 10
D21727 N21727 0 diode
R21728 N21727 N21728 10
D21728 N21728 0 diode
R21729 N21728 N21729 10
D21729 N21729 0 diode
R21730 N21729 N21730 10
D21730 N21730 0 diode
R21731 N21730 N21731 10
D21731 N21731 0 diode
R21732 N21731 N21732 10
D21732 N21732 0 diode
R21733 N21732 N21733 10
D21733 N21733 0 diode
R21734 N21733 N21734 10
D21734 N21734 0 diode
R21735 N21734 N21735 10
D21735 N21735 0 diode
R21736 N21735 N21736 10
D21736 N21736 0 diode
R21737 N21736 N21737 10
D21737 N21737 0 diode
R21738 N21737 N21738 10
D21738 N21738 0 diode
R21739 N21738 N21739 10
D21739 N21739 0 diode
R21740 N21739 N21740 10
D21740 N21740 0 diode
R21741 N21740 N21741 10
D21741 N21741 0 diode
R21742 N21741 N21742 10
D21742 N21742 0 diode
R21743 N21742 N21743 10
D21743 N21743 0 diode
R21744 N21743 N21744 10
D21744 N21744 0 diode
R21745 N21744 N21745 10
D21745 N21745 0 diode
R21746 N21745 N21746 10
D21746 N21746 0 diode
R21747 N21746 N21747 10
D21747 N21747 0 diode
R21748 N21747 N21748 10
D21748 N21748 0 diode
R21749 N21748 N21749 10
D21749 N21749 0 diode
R21750 N21749 N21750 10
D21750 N21750 0 diode
R21751 N21750 N21751 10
D21751 N21751 0 diode
R21752 N21751 N21752 10
D21752 N21752 0 diode
R21753 N21752 N21753 10
D21753 N21753 0 diode
R21754 N21753 N21754 10
D21754 N21754 0 diode
R21755 N21754 N21755 10
D21755 N21755 0 diode
R21756 N21755 N21756 10
D21756 N21756 0 diode
R21757 N21756 N21757 10
D21757 N21757 0 diode
R21758 N21757 N21758 10
D21758 N21758 0 diode
R21759 N21758 N21759 10
D21759 N21759 0 diode
R21760 N21759 N21760 10
D21760 N21760 0 diode
R21761 N21760 N21761 10
D21761 N21761 0 diode
R21762 N21761 N21762 10
D21762 N21762 0 diode
R21763 N21762 N21763 10
D21763 N21763 0 diode
R21764 N21763 N21764 10
D21764 N21764 0 diode
R21765 N21764 N21765 10
D21765 N21765 0 diode
R21766 N21765 N21766 10
D21766 N21766 0 diode
R21767 N21766 N21767 10
D21767 N21767 0 diode
R21768 N21767 N21768 10
D21768 N21768 0 diode
R21769 N21768 N21769 10
D21769 N21769 0 diode
R21770 N21769 N21770 10
D21770 N21770 0 diode
R21771 N21770 N21771 10
D21771 N21771 0 diode
R21772 N21771 N21772 10
D21772 N21772 0 diode
R21773 N21772 N21773 10
D21773 N21773 0 diode
R21774 N21773 N21774 10
D21774 N21774 0 diode
R21775 N21774 N21775 10
D21775 N21775 0 diode
R21776 N21775 N21776 10
D21776 N21776 0 diode
R21777 N21776 N21777 10
D21777 N21777 0 diode
R21778 N21777 N21778 10
D21778 N21778 0 diode
R21779 N21778 N21779 10
D21779 N21779 0 diode
R21780 N21779 N21780 10
D21780 N21780 0 diode
R21781 N21780 N21781 10
D21781 N21781 0 diode
R21782 N21781 N21782 10
D21782 N21782 0 diode
R21783 N21782 N21783 10
D21783 N21783 0 diode
R21784 N21783 N21784 10
D21784 N21784 0 diode
R21785 N21784 N21785 10
D21785 N21785 0 diode
R21786 N21785 N21786 10
D21786 N21786 0 diode
R21787 N21786 N21787 10
D21787 N21787 0 diode
R21788 N21787 N21788 10
D21788 N21788 0 diode
R21789 N21788 N21789 10
D21789 N21789 0 diode
R21790 N21789 N21790 10
D21790 N21790 0 diode
R21791 N21790 N21791 10
D21791 N21791 0 diode
R21792 N21791 N21792 10
D21792 N21792 0 diode
R21793 N21792 N21793 10
D21793 N21793 0 diode
R21794 N21793 N21794 10
D21794 N21794 0 diode
R21795 N21794 N21795 10
D21795 N21795 0 diode
R21796 N21795 N21796 10
D21796 N21796 0 diode
R21797 N21796 N21797 10
D21797 N21797 0 diode
R21798 N21797 N21798 10
D21798 N21798 0 diode
R21799 N21798 N21799 10
D21799 N21799 0 diode
R21800 N21799 N21800 10
D21800 N21800 0 diode
R21801 N21800 N21801 10
D21801 N21801 0 diode
R21802 N21801 N21802 10
D21802 N21802 0 diode
R21803 N21802 N21803 10
D21803 N21803 0 diode
R21804 N21803 N21804 10
D21804 N21804 0 diode
R21805 N21804 N21805 10
D21805 N21805 0 diode
R21806 N21805 N21806 10
D21806 N21806 0 diode
R21807 N21806 N21807 10
D21807 N21807 0 diode
R21808 N21807 N21808 10
D21808 N21808 0 diode
R21809 N21808 N21809 10
D21809 N21809 0 diode
R21810 N21809 N21810 10
D21810 N21810 0 diode
R21811 N21810 N21811 10
D21811 N21811 0 diode
R21812 N21811 N21812 10
D21812 N21812 0 diode
R21813 N21812 N21813 10
D21813 N21813 0 diode
R21814 N21813 N21814 10
D21814 N21814 0 diode
R21815 N21814 N21815 10
D21815 N21815 0 diode
R21816 N21815 N21816 10
D21816 N21816 0 diode
R21817 N21816 N21817 10
D21817 N21817 0 diode
R21818 N21817 N21818 10
D21818 N21818 0 diode
R21819 N21818 N21819 10
D21819 N21819 0 diode
R21820 N21819 N21820 10
D21820 N21820 0 diode
R21821 N21820 N21821 10
D21821 N21821 0 diode
R21822 N21821 N21822 10
D21822 N21822 0 diode
R21823 N21822 N21823 10
D21823 N21823 0 diode
R21824 N21823 N21824 10
D21824 N21824 0 diode
R21825 N21824 N21825 10
D21825 N21825 0 diode
R21826 N21825 N21826 10
D21826 N21826 0 diode
R21827 N21826 N21827 10
D21827 N21827 0 diode
R21828 N21827 N21828 10
D21828 N21828 0 diode
R21829 N21828 N21829 10
D21829 N21829 0 diode
R21830 N21829 N21830 10
D21830 N21830 0 diode
R21831 N21830 N21831 10
D21831 N21831 0 diode
R21832 N21831 N21832 10
D21832 N21832 0 diode
R21833 N21832 N21833 10
D21833 N21833 0 diode
R21834 N21833 N21834 10
D21834 N21834 0 diode
R21835 N21834 N21835 10
D21835 N21835 0 diode
R21836 N21835 N21836 10
D21836 N21836 0 diode
R21837 N21836 N21837 10
D21837 N21837 0 diode
R21838 N21837 N21838 10
D21838 N21838 0 diode
R21839 N21838 N21839 10
D21839 N21839 0 diode
R21840 N21839 N21840 10
D21840 N21840 0 diode
R21841 N21840 N21841 10
D21841 N21841 0 diode
R21842 N21841 N21842 10
D21842 N21842 0 diode
R21843 N21842 N21843 10
D21843 N21843 0 diode
R21844 N21843 N21844 10
D21844 N21844 0 diode
R21845 N21844 N21845 10
D21845 N21845 0 diode
R21846 N21845 N21846 10
D21846 N21846 0 diode
R21847 N21846 N21847 10
D21847 N21847 0 diode
R21848 N21847 N21848 10
D21848 N21848 0 diode
R21849 N21848 N21849 10
D21849 N21849 0 diode
R21850 N21849 N21850 10
D21850 N21850 0 diode
R21851 N21850 N21851 10
D21851 N21851 0 diode
R21852 N21851 N21852 10
D21852 N21852 0 diode
R21853 N21852 N21853 10
D21853 N21853 0 diode
R21854 N21853 N21854 10
D21854 N21854 0 diode
R21855 N21854 N21855 10
D21855 N21855 0 diode
R21856 N21855 N21856 10
D21856 N21856 0 diode
R21857 N21856 N21857 10
D21857 N21857 0 diode
R21858 N21857 N21858 10
D21858 N21858 0 diode
R21859 N21858 N21859 10
D21859 N21859 0 diode
R21860 N21859 N21860 10
D21860 N21860 0 diode
R21861 N21860 N21861 10
D21861 N21861 0 diode
R21862 N21861 N21862 10
D21862 N21862 0 diode
R21863 N21862 N21863 10
D21863 N21863 0 diode
R21864 N21863 N21864 10
D21864 N21864 0 diode
R21865 N21864 N21865 10
D21865 N21865 0 diode
R21866 N21865 N21866 10
D21866 N21866 0 diode
R21867 N21866 N21867 10
D21867 N21867 0 diode
R21868 N21867 N21868 10
D21868 N21868 0 diode
R21869 N21868 N21869 10
D21869 N21869 0 diode
R21870 N21869 N21870 10
D21870 N21870 0 diode
R21871 N21870 N21871 10
D21871 N21871 0 diode
R21872 N21871 N21872 10
D21872 N21872 0 diode
R21873 N21872 N21873 10
D21873 N21873 0 diode
R21874 N21873 N21874 10
D21874 N21874 0 diode
R21875 N21874 N21875 10
D21875 N21875 0 diode
R21876 N21875 N21876 10
D21876 N21876 0 diode
R21877 N21876 N21877 10
D21877 N21877 0 diode
R21878 N21877 N21878 10
D21878 N21878 0 diode
R21879 N21878 N21879 10
D21879 N21879 0 diode
R21880 N21879 N21880 10
D21880 N21880 0 diode
R21881 N21880 N21881 10
D21881 N21881 0 diode
R21882 N21881 N21882 10
D21882 N21882 0 diode
R21883 N21882 N21883 10
D21883 N21883 0 diode
R21884 N21883 N21884 10
D21884 N21884 0 diode
R21885 N21884 N21885 10
D21885 N21885 0 diode
R21886 N21885 N21886 10
D21886 N21886 0 diode
R21887 N21886 N21887 10
D21887 N21887 0 diode
R21888 N21887 N21888 10
D21888 N21888 0 diode
R21889 N21888 N21889 10
D21889 N21889 0 diode
R21890 N21889 N21890 10
D21890 N21890 0 diode
R21891 N21890 N21891 10
D21891 N21891 0 diode
R21892 N21891 N21892 10
D21892 N21892 0 diode
R21893 N21892 N21893 10
D21893 N21893 0 diode
R21894 N21893 N21894 10
D21894 N21894 0 diode
R21895 N21894 N21895 10
D21895 N21895 0 diode
R21896 N21895 N21896 10
D21896 N21896 0 diode
R21897 N21896 N21897 10
D21897 N21897 0 diode
R21898 N21897 N21898 10
D21898 N21898 0 diode
R21899 N21898 N21899 10
D21899 N21899 0 diode
R21900 N21899 N21900 10
D21900 N21900 0 diode
R21901 N21900 N21901 10
D21901 N21901 0 diode
R21902 N21901 N21902 10
D21902 N21902 0 diode
R21903 N21902 N21903 10
D21903 N21903 0 diode
R21904 N21903 N21904 10
D21904 N21904 0 diode
R21905 N21904 N21905 10
D21905 N21905 0 diode
R21906 N21905 N21906 10
D21906 N21906 0 diode
R21907 N21906 N21907 10
D21907 N21907 0 diode
R21908 N21907 N21908 10
D21908 N21908 0 diode
R21909 N21908 N21909 10
D21909 N21909 0 diode
R21910 N21909 N21910 10
D21910 N21910 0 diode
R21911 N21910 N21911 10
D21911 N21911 0 diode
R21912 N21911 N21912 10
D21912 N21912 0 diode
R21913 N21912 N21913 10
D21913 N21913 0 diode
R21914 N21913 N21914 10
D21914 N21914 0 diode
R21915 N21914 N21915 10
D21915 N21915 0 diode
R21916 N21915 N21916 10
D21916 N21916 0 diode
R21917 N21916 N21917 10
D21917 N21917 0 diode
R21918 N21917 N21918 10
D21918 N21918 0 diode
R21919 N21918 N21919 10
D21919 N21919 0 diode
R21920 N21919 N21920 10
D21920 N21920 0 diode
R21921 N21920 N21921 10
D21921 N21921 0 diode
R21922 N21921 N21922 10
D21922 N21922 0 diode
R21923 N21922 N21923 10
D21923 N21923 0 diode
R21924 N21923 N21924 10
D21924 N21924 0 diode
R21925 N21924 N21925 10
D21925 N21925 0 diode
R21926 N21925 N21926 10
D21926 N21926 0 diode
R21927 N21926 N21927 10
D21927 N21927 0 diode
R21928 N21927 N21928 10
D21928 N21928 0 diode
R21929 N21928 N21929 10
D21929 N21929 0 diode
R21930 N21929 N21930 10
D21930 N21930 0 diode
R21931 N21930 N21931 10
D21931 N21931 0 diode
R21932 N21931 N21932 10
D21932 N21932 0 diode
R21933 N21932 N21933 10
D21933 N21933 0 diode
R21934 N21933 N21934 10
D21934 N21934 0 diode
R21935 N21934 N21935 10
D21935 N21935 0 diode
R21936 N21935 N21936 10
D21936 N21936 0 diode
R21937 N21936 N21937 10
D21937 N21937 0 diode
R21938 N21937 N21938 10
D21938 N21938 0 diode
R21939 N21938 N21939 10
D21939 N21939 0 diode
R21940 N21939 N21940 10
D21940 N21940 0 diode
R21941 N21940 N21941 10
D21941 N21941 0 diode
R21942 N21941 N21942 10
D21942 N21942 0 diode
R21943 N21942 N21943 10
D21943 N21943 0 diode
R21944 N21943 N21944 10
D21944 N21944 0 diode
R21945 N21944 N21945 10
D21945 N21945 0 diode
R21946 N21945 N21946 10
D21946 N21946 0 diode
R21947 N21946 N21947 10
D21947 N21947 0 diode
R21948 N21947 N21948 10
D21948 N21948 0 diode
R21949 N21948 N21949 10
D21949 N21949 0 diode
R21950 N21949 N21950 10
D21950 N21950 0 diode
R21951 N21950 N21951 10
D21951 N21951 0 diode
R21952 N21951 N21952 10
D21952 N21952 0 diode
R21953 N21952 N21953 10
D21953 N21953 0 diode
R21954 N21953 N21954 10
D21954 N21954 0 diode
R21955 N21954 N21955 10
D21955 N21955 0 diode
R21956 N21955 N21956 10
D21956 N21956 0 diode
R21957 N21956 N21957 10
D21957 N21957 0 diode
R21958 N21957 N21958 10
D21958 N21958 0 diode
R21959 N21958 N21959 10
D21959 N21959 0 diode
R21960 N21959 N21960 10
D21960 N21960 0 diode
R21961 N21960 N21961 10
D21961 N21961 0 diode
R21962 N21961 N21962 10
D21962 N21962 0 diode
R21963 N21962 N21963 10
D21963 N21963 0 diode
R21964 N21963 N21964 10
D21964 N21964 0 diode
R21965 N21964 N21965 10
D21965 N21965 0 diode
R21966 N21965 N21966 10
D21966 N21966 0 diode
R21967 N21966 N21967 10
D21967 N21967 0 diode
R21968 N21967 N21968 10
D21968 N21968 0 diode
R21969 N21968 N21969 10
D21969 N21969 0 diode
R21970 N21969 N21970 10
D21970 N21970 0 diode
R21971 N21970 N21971 10
D21971 N21971 0 diode
R21972 N21971 N21972 10
D21972 N21972 0 diode
R21973 N21972 N21973 10
D21973 N21973 0 diode
R21974 N21973 N21974 10
D21974 N21974 0 diode
R21975 N21974 N21975 10
D21975 N21975 0 diode
R21976 N21975 N21976 10
D21976 N21976 0 diode
R21977 N21976 N21977 10
D21977 N21977 0 diode
R21978 N21977 N21978 10
D21978 N21978 0 diode
R21979 N21978 N21979 10
D21979 N21979 0 diode
R21980 N21979 N21980 10
D21980 N21980 0 diode
R21981 N21980 N21981 10
D21981 N21981 0 diode
R21982 N21981 N21982 10
D21982 N21982 0 diode
R21983 N21982 N21983 10
D21983 N21983 0 diode
R21984 N21983 N21984 10
D21984 N21984 0 diode
R21985 N21984 N21985 10
D21985 N21985 0 diode
R21986 N21985 N21986 10
D21986 N21986 0 diode
R21987 N21986 N21987 10
D21987 N21987 0 diode
R21988 N21987 N21988 10
D21988 N21988 0 diode
R21989 N21988 N21989 10
D21989 N21989 0 diode
R21990 N21989 N21990 10
D21990 N21990 0 diode
R21991 N21990 N21991 10
D21991 N21991 0 diode
R21992 N21991 N21992 10
D21992 N21992 0 diode
R21993 N21992 N21993 10
D21993 N21993 0 diode
R21994 N21993 N21994 10
D21994 N21994 0 diode
R21995 N21994 N21995 10
D21995 N21995 0 diode
R21996 N21995 N21996 10
D21996 N21996 0 diode
R21997 N21996 N21997 10
D21997 N21997 0 diode
R21998 N21997 N21998 10
D21998 N21998 0 diode
R21999 N21998 N21999 10
D21999 N21999 0 diode
R22000 N21999 N22000 10
D22000 N22000 0 diode
R22001 N22000 N22001 10
D22001 N22001 0 diode
R22002 N22001 N22002 10
D22002 N22002 0 diode
R22003 N22002 N22003 10
D22003 N22003 0 diode
R22004 N22003 N22004 10
D22004 N22004 0 diode
R22005 N22004 N22005 10
D22005 N22005 0 diode
R22006 N22005 N22006 10
D22006 N22006 0 diode
R22007 N22006 N22007 10
D22007 N22007 0 diode
R22008 N22007 N22008 10
D22008 N22008 0 diode
R22009 N22008 N22009 10
D22009 N22009 0 diode
R22010 N22009 N22010 10
D22010 N22010 0 diode
R22011 N22010 N22011 10
D22011 N22011 0 diode
R22012 N22011 N22012 10
D22012 N22012 0 diode
R22013 N22012 N22013 10
D22013 N22013 0 diode
R22014 N22013 N22014 10
D22014 N22014 0 diode
R22015 N22014 N22015 10
D22015 N22015 0 diode
R22016 N22015 N22016 10
D22016 N22016 0 diode
R22017 N22016 N22017 10
D22017 N22017 0 diode
R22018 N22017 N22018 10
D22018 N22018 0 diode
R22019 N22018 N22019 10
D22019 N22019 0 diode
R22020 N22019 N22020 10
D22020 N22020 0 diode
R22021 N22020 N22021 10
D22021 N22021 0 diode
R22022 N22021 N22022 10
D22022 N22022 0 diode
R22023 N22022 N22023 10
D22023 N22023 0 diode
R22024 N22023 N22024 10
D22024 N22024 0 diode
R22025 N22024 N22025 10
D22025 N22025 0 diode
R22026 N22025 N22026 10
D22026 N22026 0 diode
R22027 N22026 N22027 10
D22027 N22027 0 diode
R22028 N22027 N22028 10
D22028 N22028 0 diode
R22029 N22028 N22029 10
D22029 N22029 0 diode
R22030 N22029 N22030 10
D22030 N22030 0 diode
R22031 N22030 N22031 10
D22031 N22031 0 diode
R22032 N22031 N22032 10
D22032 N22032 0 diode
R22033 N22032 N22033 10
D22033 N22033 0 diode
R22034 N22033 N22034 10
D22034 N22034 0 diode
R22035 N22034 N22035 10
D22035 N22035 0 diode
R22036 N22035 N22036 10
D22036 N22036 0 diode
R22037 N22036 N22037 10
D22037 N22037 0 diode
R22038 N22037 N22038 10
D22038 N22038 0 diode
R22039 N22038 N22039 10
D22039 N22039 0 diode
R22040 N22039 N22040 10
D22040 N22040 0 diode
R22041 N22040 N22041 10
D22041 N22041 0 diode
R22042 N22041 N22042 10
D22042 N22042 0 diode
R22043 N22042 N22043 10
D22043 N22043 0 diode
R22044 N22043 N22044 10
D22044 N22044 0 diode
R22045 N22044 N22045 10
D22045 N22045 0 diode
R22046 N22045 N22046 10
D22046 N22046 0 diode
R22047 N22046 N22047 10
D22047 N22047 0 diode
R22048 N22047 N22048 10
D22048 N22048 0 diode
R22049 N22048 N22049 10
D22049 N22049 0 diode
R22050 N22049 N22050 10
D22050 N22050 0 diode
R22051 N22050 N22051 10
D22051 N22051 0 diode
R22052 N22051 N22052 10
D22052 N22052 0 diode
R22053 N22052 N22053 10
D22053 N22053 0 diode
R22054 N22053 N22054 10
D22054 N22054 0 diode
R22055 N22054 N22055 10
D22055 N22055 0 diode
R22056 N22055 N22056 10
D22056 N22056 0 diode
R22057 N22056 N22057 10
D22057 N22057 0 diode
R22058 N22057 N22058 10
D22058 N22058 0 diode
R22059 N22058 N22059 10
D22059 N22059 0 diode
R22060 N22059 N22060 10
D22060 N22060 0 diode
R22061 N22060 N22061 10
D22061 N22061 0 diode
R22062 N22061 N22062 10
D22062 N22062 0 diode
R22063 N22062 N22063 10
D22063 N22063 0 diode
R22064 N22063 N22064 10
D22064 N22064 0 diode
R22065 N22064 N22065 10
D22065 N22065 0 diode
R22066 N22065 N22066 10
D22066 N22066 0 diode
R22067 N22066 N22067 10
D22067 N22067 0 diode
R22068 N22067 N22068 10
D22068 N22068 0 diode
R22069 N22068 N22069 10
D22069 N22069 0 diode
R22070 N22069 N22070 10
D22070 N22070 0 diode
R22071 N22070 N22071 10
D22071 N22071 0 diode
R22072 N22071 N22072 10
D22072 N22072 0 diode
R22073 N22072 N22073 10
D22073 N22073 0 diode
R22074 N22073 N22074 10
D22074 N22074 0 diode
R22075 N22074 N22075 10
D22075 N22075 0 diode
R22076 N22075 N22076 10
D22076 N22076 0 diode
R22077 N22076 N22077 10
D22077 N22077 0 diode
R22078 N22077 N22078 10
D22078 N22078 0 diode
R22079 N22078 N22079 10
D22079 N22079 0 diode
R22080 N22079 N22080 10
D22080 N22080 0 diode
R22081 N22080 N22081 10
D22081 N22081 0 diode
R22082 N22081 N22082 10
D22082 N22082 0 diode
R22083 N22082 N22083 10
D22083 N22083 0 diode
R22084 N22083 N22084 10
D22084 N22084 0 diode
R22085 N22084 N22085 10
D22085 N22085 0 diode
R22086 N22085 N22086 10
D22086 N22086 0 diode
R22087 N22086 N22087 10
D22087 N22087 0 diode
R22088 N22087 N22088 10
D22088 N22088 0 diode
R22089 N22088 N22089 10
D22089 N22089 0 diode
R22090 N22089 N22090 10
D22090 N22090 0 diode
R22091 N22090 N22091 10
D22091 N22091 0 diode
R22092 N22091 N22092 10
D22092 N22092 0 diode
R22093 N22092 N22093 10
D22093 N22093 0 diode
R22094 N22093 N22094 10
D22094 N22094 0 diode
R22095 N22094 N22095 10
D22095 N22095 0 diode
R22096 N22095 N22096 10
D22096 N22096 0 diode
R22097 N22096 N22097 10
D22097 N22097 0 diode
R22098 N22097 N22098 10
D22098 N22098 0 diode
R22099 N22098 N22099 10
D22099 N22099 0 diode
R22100 N22099 N22100 10
D22100 N22100 0 diode
R22101 N22100 N22101 10
D22101 N22101 0 diode
R22102 N22101 N22102 10
D22102 N22102 0 diode
R22103 N22102 N22103 10
D22103 N22103 0 diode
R22104 N22103 N22104 10
D22104 N22104 0 diode
R22105 N22104 N22105 10
D22105 N22105 0 diode
R22106 N22105 N22106 10
D22106 N22106 0 diode
R22107 N22106 N22107 10
D22107 N22107 0 diode
R22108 N22107 N22108 10
D22108 N22108 0 diode
R22109 N22108 N22109 10
D22109 N22109 0 diode
R22110 N22109 N22110 10
D22110 N22110 0 diode
R22111 N22110 N22111 10
D22111 N22111 0 diode
R22112 N22111 N22112 10
D22112 N22112 0 diode
R22113 N22112 N22113 10
D22113 N22113 0 diode
R22114 N22113 N22114 10
D22114 N22114 0 diode
R22115 N22114 N22115 10
D22115 N22115 0 diode
R22116 N22115 N22116 10
D22116 N22116 0 diode
R22117 N22116 N22117 10
D22117 N22117 0 diode
R22118 N22117 N22118 10
D22118 N22118 0 diode
R22119 N22118 N22119 10
D22119 N22119 0 diode
R22120 N22119 N22120 10
D22120 N22120 0 diode
R22121 N22120 N22121 10
D22121 N22121 0 diode
R22122 N22121 N22122 10
D22122 N22122 0 diode
R22123 N22122 N22123 10
D22123 N22123 0 diode
R22124 N22123 N22124 10
D22124 N22124 0 diode
R22125 N22124 N22125 10
D22125 N22125 0 diode
R22126 N22125 N22126 10
D22126 N22126 0 diode
R22127 N22126 N22127 10
D22127 N22127 0 diode
R22128 N22127 N22128 10
D22128 N22128 0 diode
R22129 N22128 N22129 10
D22129 N22129 0 diode
R22130 N22129 N22130 10
D22130 N22130 0 diode
R22131 N22130 N22131 10
D22131 N22131 0 diode
R22132 N22131 N22132 10
D22132 N22132 0 diode
R22133 N22132 N22133 10
D22133 N22133 0 diode
R22134 N22133 N22134 10
D22134 N22134 0 diode
R22135 N22134 N22135 10
D22135 N22135 0 diode
R22136 N22135 N22136 10
D22136 N22136 0 diode
R22137 N22136 N22137 10
D22137 N22137 0 diode
R22138 N22137 N22138 10
D22138 N22138 0 diode
R22139 N22138 N22139 10
D22139 N22139 0 diode
R22140 N22139 N22140 10
D22140 N22140 0 diode
R22141 N22140 N22141 10
D22141 N22141 0 diode
R22142 N22141 N22142 10
D22142 N22142 0 diode
R22143 N22142 N22143 10
D22143 N22143 0 diode
R22144 N22143 N22144 10
D22144 N22144 0 diode
R22145 N22144 N22145 10
D22145 N22145 0 diode
R22146 N22145 N22146 10
D22146 N22146 0 diode
R22147 N22146 N22147 10
D22147 N22147 0 diode
R22148 N22147 N22148 10
D22148 N22148 0 diode
R22149 N22148 N22149 10
D22149 N22149 0 diode
R22150 N22149 N22150 10
D22150 N22150 0 diode
R22151 N22150 N22151 10
D22151 N22151 0 diode
R22152 N22151 N22152 10
D22152 N22152 0 diode
R22153 N22152 N22153 10
D22153 N22153 0 diode
R22154 N22153 N22154 10
D22154 N22154 0 diode
R22155 N22154 N22155 10
D22155 N22155 0 diode
R22156 N22155 N22156 10
D22156 N22156 0 diode
R22157 N22156 N22157 10
D22157 N22157 0 diode
R22158 N22157 N22158 10
D22158 N22158 0 diode
R22159 N22158 N22159 10
D22159 N22159 0 diode
R22160 N22159 N22160 10
D22160 N22160 0 diode
R22161 N22160 N22161 10
D22161 N22161 0 diode
R22162 N22161 N22162 10
D22162 N22162 0 diode
R22163 N22162 N22163 10
D22163 N22163 0 diode
R22164 N22163 N22164 10
D22164 N22164 0 diode
R22165 N22164 N22165 10
D22165 N22165 0 diode
R22166 N22165 N22166 10
D22166 N22166 0 diode
R22167 N22166 N22167 10
D22167 N22167 0 diode
R22168 N22167 N22168 10
D22168 N22168 0 diode
R22169 N22168 N22169 10
D22169 N22169 0 diode
R22170 N22169 N22170 10
D22170 N22170 0 diode
R22171 N22170 N22171 10
D22171 N22171 0 diode
R22172 N22171 N22172 10
D22172 N22172 0 diode
R22173 N22172 N22173 10
D22173 N22173 0 diode
R22174 N22173 N22174 10
D22174 N22174 0 diode
R22175 N22174 N22175 10
D22175 N22175 0 diode
R22176 N22175 N22176 10
D22176 N22176 0 diode
R22177 N22176 N22177 10
D22177 N22177 0 diode
R22178 N22177 N22178 10
D22178 N22178 0 diode
R22179 N22178 N22179 10
D22179 N22179 0 diode
R22180 N22179 N22180 10
D22180 N22180 0 diode
R22181 N22180 N22181 10
D22181 N22181 0 diode
R22182 N22181 N22182 10
D22182 N22182 0 diode
R22183 N22182 N22183 10
D22183 N22183 0 diode
R22184 N22183 N22184 10
D22184 N22184 0 diode
R22185 N22184 N22185 10
D22185 N22185 0 diode
R22186 N22185 N22186 10
D22186 N22186 0 diode
R22187 N22186 N22187 10
D22187 N22187 0 diode
R22188 N22187 N22188 10
D22188 N22188 0 diode
R22189 N22188 N22189 10
D22189 N22189 0 diode
R22190 N22189 N22190 10
D22190 N22190 0 diode
R22191 N22190 N22191 10
D22191 N22191 0 diode
R22192 N22191 N22192 10
D22192 N22192 0 diode
R22193 N22192 N22193 10
D22193 N22193 0 diode
R22194 N22193 N22194 10
D22194 N22194 0 diode
R22195 N22194 N22195 10
D22195 N22195 0 diode
R22196 N22195 N22196 10
D22196 N22196 0 diode
R22197 N22196 N22197 10
D22197 N22197 0 diode
R22198 N22197 N22198 10
D22198 N22198 0 diode
R22199 N22198 N22199 10
D22199 N22199 0 diode
R22200 N22199 N22200 10
D22200 N22200 0 diode
R22201 N22200 N22201 10
D22201 N22201 0 diode
R22202 N22201 N22202 10
D22202 N22202 0 diode
R22203 N22202 N22203 10
D22203 N22203 0 diode
R22204 N22203 N22204 10
D22204 N22204 0 diode
R22205 N22204 N22205 10
D22205 N22205 0 diode
R22206 N22205 N22206 10
D22206 N22206 0 diode
R22207 N22206 N22207 10
D22207 N22207 0 diode
R22208 N22207 N22208 10
D22208 N22208 0 diode
R22209 N22208 N22209 10
D22209 N22209 0 diode
R22210 N22209 N22210 10
D22210 N22210 0 diode
R22211 N22210 N22211 10
D22211 N22211 0 diode
R22212 N22211 N22212 10
D22212 N22212 0 diode
R22213 N22212 N22213 10
D22213 N22213 0 diode
R22214 N22213 N22214 10
D22214 N22214 0 diode
R22215 N22214 N22215 10
D22215 N22215 0 diode
R22216 N22215 N22216 10
D22216 N22216 0 diode
R22217 N22216 N22217 10
D22217 N22217 0 diode
R22218 N22217 N22218 10
D22218 N22218 0 diode
R22219 N22218 N22219 10
D22219 N22219 0 diode
R22220 N22219 N22220 10
D22220 N22220 0 diode
R22221 N22220 N22221 10
D22221 N22221 0 diode
R22222 N22221 N22222 10
D22222 N22222 0 diode
R22223 N22222 N22223 10
D22223 N22223 0 diode
R22224 N22223 N22224 10
D22224 N22224 0 diode
R22225 N22224 N22225 10
D22225 N22225 0 diode
R22226 N22225 N22226 10
D22226 N22226 0 diode
R22227 N22226 N22227 10
D22227 N22227 0 diode
R22228 N22227 N22228 10
D22228 N22228 0 diode
R22229 N22228 N22229 10
D22229 N22229 0 diode
R22230 N22229 N22230 10
D22230 N22230 0 diode
R22231 N22230 N22231 10
D22231 N22231 0 diode
R22232 N22231 N22232 10
D22232 N22232 0 diode
R22233 N22232 N22233 10
D22233 N22233 0 diode
R22234 N22233 N22234 10
D22234 N22234 0 diode
R22235 N22234 N22235 10
D22235 N22235 0 diode
R22236 N22235 N22236 10
D22236 N22236 0 diode
R22237 N22236 N22237 10
D22237 N22237 0 diode
R22238 N22237 N22238 10
D22238 N22238 0 diode
R22239 N22238 N22239 10
D22239 N22239 0 diode
R22240 N22239 N22240 10
D22240 N22240 0 diode
R22241 N22240 N22241 10
D22241 N22241 0 diode
R22242 N22241 N22242 10
D22242 N22242 0 diode
R22243 N22242 N22243 10
D22243 N22243 0 diode
R22244 N22243 N22244 10
D22244 N22244 0 diode
R22245 N22244 N22245 10
D22245 N22245 0 diode
R22246 N22245 N22246 10
D22246 N22246 0 diode
R22247 N22246 N22247 10
D22247 N22247 0 diode
R22248 N22247 N22248 10
D22248 N22248 0 diode
R22249 N22248 N22249 10
D22249 N22249 0 diode
R22250 N22249 N22250 10
D22250 N22250 0 diode
R22251 N22250 N22251 10
D22251 N22251 0 diode
R22252 N22251 N22252 10
D22252 N22252 0 diode
R22253 N22252 N22253 10
D22253 N22253 0 diode
R22254 N22253 N22254 10
D22254 N22254 0 diode
R22255 N22254 N22255 10
D22255 N22255 0 diode
R22256 N22255 N22256 10
D22256 N22256 0 diode
R22257 N22256 N22257 10
D22257 N22257 0 diode
R22258 N22257 N22258 10
D22258 N22258 0 diode
R22259 N22258 N22259 10
D22259 N22259 0 diode
R22260 N22259 N22260 10
D22260 N22260 0 diode
R22261 N22260 N22261 10
D22261 N22261 0 diode
R22262 N22261 N22262 10
D22262 N22262 0 diode
R22263 N22262 N22263 10
D22263 N22263 0 diode
R22264 N22263 N22264 10
D22264 N22264 0 diode
R22265 N22264 N22265 10
D22265 N22265 0 diode
R22266 N22265 N22266 10
D22266 N22266 0 diode
R22267 N22266 N22267 10
D22267 N22267 0 diode
R22268 N22267 N22268 10
D22268 N22268 0 diode
R22269 N22268 N22269 10
D22269 N22269 0 diode
R22270 N22269 N22270 10
D22270 N22270 0 diode
R22271 N22270 N22271 10
D22271 N22271 0 diode
R22272 N22271 N22272 10
D22272 N22272 0 diode
R22273 N22272 N22273 10
D22273 N22273 0 diode
R22274 N22273 N22274 10
D22274 N22274 0 diode
R22275 N22274 N22275 10
D22275 N22275 0 diode
R22276 N22275 N22276 10
D22276 N22276 0 diode
R22277 N22276 N22277 10
D22277 N22277 0 diode
R22278 N22277 N22278 10
D22278 N22278 0 diode
R22279 N22278 N22279 10
D22279 N22279 0 diode
R22280 N22279 N22280 10
D22280 N22280 0 diode
R22281 N22280 N22281 10
D22281 N22281 0 diode
R22282 N22281 N22282 10
D22282 N22282 0 diode
R22283 N22282 N22283 10
D22283 N22283 0 diode
R22284 N22283 N22284 10
D22284 N22284 0 diode
R22285 N22284 N22285 10
D22285 N22285 0 diode
R22286 N22285 N22286 10
D22286 N22286 0 diode
R22287 N22286 N22287 10
D22287 N22287 0 diode
R22288 N22287 N22288 10
D22288 N22288 0 diode
R22289 N22288 N22289 10
D22289 N22289 0 diode
R22290 N22289 N22290 10
D22290 N22290 0 diode
R22291 N22290 N22291 10
D22291 N22291 0 diode
R22292 N22291 N22292 10
D22292 N22292 0 diode
R22293 N22292 N22293 10
D22293 N22293 0 diode
R22294 N22293 N22294 10
D22294 N22294 0 diode
R22295 N22294 N22295 10
D22295 N22295 0 diode
R22296 N22295 N22296 10
D22296 N22296 0 diode
R22297 N22296 N22297 10
D22297 N22297 0 diode
R22298 N22297 N22298 10
D22298 N22298 0 diode
R22299 N22298 N22299 10
D22299 N22299 0 diode
R22300 N22299 N22300 10
D22300 N22300 0 diode
R22301 N22300 N22301 10
D22301 N22301 0 diode
R22302 N22301 N22302 10
D22302 N22302 0 diode
R22303 N22302 N22303 10
D22303 N22303 0 diode
R22304 N22303 N22304 10
D22304 N22304 0 diode
R22305 N22304 N22305 10
D22305 N22305 0 diode
R22306 N22305 N22306 10
D22306 N22306 0 diode
R22307 N22306 N22307 10
D22307 N22307 0 diode
R22308 N22307 N22308 10
D22308 N22308 0 diode
R22309 N22308 N22309 10
D22309 N22309 0 diode
R22310 N22309 N22310 10
D22310 N22310 0 diode
R22311 N22310 N22311 10
D22311 N22311 0 diode
R22312 N22311 N22312 10
D22312 N22312 0 diode
R22313 N22312 N22313 10
D22313 N22313 0 diode
R22314 N22313 N22314 10
D22314 N22314 0 diode
R22315 N22314 N22315 10
D22315 N22315 0 diode
R22316 N22315 N22316 10
D22316 N22316 0 diode
R22317 N22316 N22317 10
D22317 N22317 0 diode
R22318 N22317 N22318 10
D22318 N22318 0 diode
R22319 N22318 N22319 10
D22319 N22319 0 diode
R22320 N22319 N22320 10
D22320 N22320 0 diode
R22321 N22320 N22321 10
D22321 N22321 0 diode
R22322 N22321 N22322 10
D22322 N22322 0 diode
R22323 N22322 N22323 10
D22323 N22323 0 diode
R22324 N22323 N22324 10
D22324 N22324 0 diode
R22325 N22324 N22325 10
D22325 N22325 0 diode
R22326 N22325 N22326 10
D22326 N22326 0 diode
R22327 N22326 N22327 10
D22327 N22327 0 diode
R22328 N22327 N22328 10
D22328 N22328 0 diode
R22329 N22328 N22329 10
D22329 N22329 0 diode
R22330 N22329 N22330 10
D22330 N22330 0 diode
R22331 N22330 N22331 10
D22331 N22331 0 diode
R22332 N22331 N22332 10
D22332 N22332 0 diode
R22333 N22332 N22333 10
D22333 N22333 0 diode
R22334 N22333 N22334 10
D22334 N22334 0 diode
R22335 N22334 N22335 10
D22335 N22335 0 diode
R22336 N22335 N22336 10
D22336 N22336 0 diode
R22337 N22336 N22337 10
D22337 N22337 0 diode
R22338 N22337 N22338 10
D22338 N22338 0 diode
R22339 N22338 N22339 10
D22339 N22339 0 diode
R22340 N22339 N22340 10
D22340 N22340 0 diode
R22341 N22340 N22341 10
D22341 N22341 0 diode
R22342 N22341 N22342 10
D22342 N22342 0 diode
R22343 N22342 N22343 10
D22343 N22343 0 diode
R22344 N22343 N22344 10
D22344 N22344 0 diode
R22345 N22344 N22345 10
D22345 N22345 0 diode
R22346 N22345 N22346 10
D22346 N22346 0 diode
R22347 N22346 N22347 10
D22347 N22347 0 diode
R22348 N22347 N22348 10
D22348 N22348 0 diode
R22349 N22348 N22349 10
D22349 N22349 0 diode
R22350 N22349 N22350 10
D22350 N22350 0 diode
R22351 N22350 N22351 10
D22351 N22351 0 diode
R22352 N22351 N22352 10
D22352 N22352 0 diode
R22353 N22352 N22353 10
D22353 N22353 0 diode
R22354 N22353 N22354 10
D22354 N22354 0 diode
R22355 N22354 N22355 10
D22355 N22355 0 diode
R22356 N22355 N22356 10
D22356 N22356 0 diode
R22357 N22356 N22357 10
D22357 N22357 0 diode
R22358 N22357 N22358 10
D22358 N22358 0 diode
R22359 N22358 N22359 10
D22359 N22359 0 diode
R22360 N22359 N22360 10
D22360 N22360 0 diode
R22361 N22360 N22361 10
D22361 N22361 0 diode
R22362 N22361 N22362 10
D22362 N22362 0 diode
R22363 N22362 N22363 10
D22363 N22363 0 diode
R22364 N22363 N22364 10
D22364 N22364 0 diode
R22365 N22364 N22365 10
D22365 N22365 0 diode
R22366 N22365 N22366 10
D22366 N22366 0 diode
R22367 N22366 N22367 10
D22367 N22367 0 diode
R22368 N22367 N22368 10
D22368 N22368 0 diode
R22369 N22368 N22369 10
D22369 N22369 0 diode
R22370 N22369 N22370 10
D22370 N22370 0 diode
R22371 N22370 N22371 10
D22371 N22371 0 diode
R22372 N22371 N22372 10
D22372 N22372 0 diode
R22373 N22372 N22373 10
D22373 N22373 0 diode
R22374 N22373 N22374 10
D22374 N22374 0 diode
R22375 N22374 N22375 10
D22375 N22375 0 diode
R22376 N22375 N22376 10
D22376 N22376 0 diode
R22377 N22376 N22377 10
D22377 N22377 0 diode
R22378 N22377 N22378 10
D22378 N22378 0 diode
R22379 N22378 N22379 10
D22379 N22379 0 diode
R22380 N22379 N22380 10
D22380 N22380 0 diode
R22381 N22380 N22381 10
D22381 N22381 0 diode
R22382 N22381 N22382 10
D22382 N22382 0 diode
R22383 N22382 N22383 10
D22383 N22383 0 diode
R22384 N22383 N22384 10
D22384 N22384 0 diode
R22385 N22384 N22385 10
D22385 N22385 0 diode
R22386 N22385 N22386 10
D22386 N22386 0 diode
R22387 N22386 N22387 10
D22387 N22387 0 diode
R22388 N22387 N22388 10
D22388 N22388 0 diode
R22389 N22388 N22389 10
D22389 N22389 0 diode
R22390 N22389 N22390 10
D22390 N22390 0 diode
R22391 N22390 N22391 10
D22391 N22391 0 diode
R22392 N22391 N22392 10
D22392 N22392 0 diode
R22393 N22392 N22393 10
D22393 N22393 0 diode
R22394 N22393 N22394 10
D22394 N22394 0 diode
R22395 N22394 N22395 10
D22395 N22395 0 diode
R22396 N22395 N22396 10
D22396 N22396 0 diode
R22397 N22396 N22397 10
D22397 N22397 0 diode
R22398 N22397 N22398 10
D22398 N22398 0 diode
R22399 N22398 N22399 10
D22399 N22399 0 diode
R22400 N22399 N22400 10
D22400 N22400 0 diode
R22401 N22400 N22401 10
D22401 N22401 0 diode
R22402 N22401 N22402 10
D22402 N22402 0 diode
R22403 N22402 N22403 10
D22403 N22403 0 diode
R22404 N22403 N22404 10
D22404 N22404 0 diode
R22405 N22404 N22405 10
D22405 N22405 0 diode
R22406 N22405 N22406 10
D22406 N22406 0 diode
R22407 N22406 N22407 10
D22407 N22407 0 diode
R22408 N22407 N22408 10
D22408 N22408 0 diode
R22409 N22408 N22409 10
D22409 N22409 0 diode
R22410 N22409 N22410 10
D22410 N22410 0 diode
R22411 N22410 N22411 10
D22411 N22411 0 diode
R22412 N22411 N22412 10
D22412 N22412 0 diode
R22413 N22412 N22413 10
D22413 N22413 0 diode
R22414 N22413 N22414 10
D22414 N22414 0 diode
R22415 N22414 N22415 10
D22415 N22415 0 diode
R22416 N22415 N22416 10
D22416 N22416 0 diode
R22417 N22416 N22417 10
D22417 N22417 0 diode
R22418 N22417 N22418 10
D22418 N22418 0 diode
R22419 N22418 N22419 10
D22419 N22419 0 diode
R22420 N22419 N22420 10
D22420 N22420 0 diode
R22421 N22420 N22421 10
D22421 N22421 0 diode
R22422 N22421 N22422 10
D22422 N22422 0 diode
R22423 N22422 N22423 10
D22423 N22423 0 diode
R22424 N22423 N22424 10
D22424 N22424 0 diode
R22425 N22424 N22425 10
D22425 N22425 0 diode
R22426 N22425 N22426 10
D22426 N22426 0 diode
R22427 N22426 N22427 10
D22427 N22427 0 diode
R22428 N22427 N22428 10
D22428 N22428 0 diode
R22429 N22428 N22429 10
D22429 N22429 0 diode
R22430 N22429 N22430 10
D22430 N22430 0 diode
R22431 N22430 N22431 10
D22431 N22431 0 diode
R22432 N22431 N22432 10
D22432 N22432 0 diode
R22433 N22432 N22433 10
D22433 N22433 0 diode
R22434 N22433 N22434 10
D22434 N22434 0 diode
R22435 N22434 N22435 10
D22435 N22435 0 diode
R22436 N22435 N22436 10
D22436 N22436 0 diode
R22437 N22436 N22437 10
D22437 N22437 0 diode
R22438 N22437 N22438 10
D22438 N22438 0 diode
R22439 N22438 N22439 10
D22439 N22439 0 diode
R22440 N22439 N22440 10
D22440 N22440 0 diode
R22441 N22440 N22441 10
D22441 N22441 0 diode
R22442 N22441 N22442 10
D22442 N22442 0 diode
R22443 N22442 N22443 10
D22443 N22443 0 diode
R22444 N22443 N22444 10
D22444 N22444 0 diode
R22445 N22444 N22445 10
D22445 N22445 0 diode
R22446 N22445 N22446 10
D22446 N22446 0 diode
R22447 N22446 N22447 10
D22447 N22447 0 diode
R22448 N22447 N22448 10
D22448 N22448 0 diode
R22449 N22448 N22449 10
D22449 N22449 0 diode
R22450 N22449 N22450 10
D22450 N22450 0 diode
R22451 N22450 N22451 10
D22451 N22451 0 diode
R22452 N22451 N22452 10
D22452 N22452 0 diode
R22453 N22452 N22453 10
D22453 N22453 0 diode
R22454 N22453 N22454 10
D22454 N22454 0 diode
R22455 N22454 N22455 10
D22455 N22455 0 diode
R22456 N22455 N22456 10
D22456 N22456 0 diode
R22457 N22456 N22457 10
D22457 N22457 0 diode
R22458 N22457 N22458 10
D22458 N22458 0 diode
R22459 N22458 N22459 10
D22459 N22459 0 diode
R22460 N22459 N22460 10
D22460 N22460 0 diode
R22461 N22460 N22461 10
D22461 N22461 0 diode
R22462 N22461 N22462 10
D22462 N22462 0 diode
R22463 N22462 N22463 10
D22463 N22463 0 diode
R22464 N22463 N22464 10
D22464 N22464 0 diode
R22465 N22464 N22465 10
D22465 N22465 0 diode
R22466 N22465 N22466 10
D22466 N22466 0 diode
R22467 N22466 N22467 10
D22467 N22467 0 diode
R22468 N22467 N22468 10
D22468 N22468 0 diode
R22469 N22468 N22469 10
D22469 N22469 0 diode
R22470 N22469 N22470 10
D22470 N22470 0 diode
R22471 N22470 N22471 10
D22471 N22471 0 diode
R22472 N22471 N22472 10
D22472 N22472 0 diode
R22473 N22472 N22473 10
D22473 N22473 0 diode
R22474 N22473 N22474 10
D22474 N22474 0 diode
R22475 N22474 N22475 10
D22475 N22475 0 diode
R22476 N22475 N22476 10
D22476 N22476 0 diode
R22477 N22476 N22477 10
D22477 N22477 0 diode
R22478 N22477 N22478 10
D22478 N22478 0 diode
R22479 N22478 N22479 10
D22479 N22479 0 diode
R22480 N22479 N22480 10
D22480 N22480 0 diode
R22481 N22480 N22481 10
D22481 N22481 0 diode
R22482 N22481 N22482 10
D22482 N22482 0 diode
R22483 N22482 N22483 10
D22483 N22483 0 diode
R22484 N22483 N22484 10
D22484 N22484 0 diode
R22485 N22484 N22485 10
D22485 N22485 0 diode
R22486 N22485 N22486 10
D22486 N22486 0 diode
R22487 N22486 N22487 10
D22487 N22487 0 diode
R22488 N22487 N22488 10
D22488 N22488 0 diode
R22489 N22488 N22489 10
D22489 N22489 0 diode
R22490 N22489 N22490 10
D22490 N22490 0 diode
R22491 N22490 N22491 10
D22491 N22491 0 diode
R22492 N22491 N22492 10
D22492 N22492 0 diode
R22493 N22492 N22493 10
D22493 N22493 0 diode
R22494 N22493 N22494 10
D22494 N22494 0 diode
R22495 N22494 N22495 10
D22495 N22495 0 diode
R22496 N22495 N22496 10
D22496 N22496 0 diode
R22497 N22496 N22497 10
D22497 N22497 0 diode
R22498 N22497 N22498 10
D22498 N22498 0 diode
R22499 N22498 N22499 10
D22499 N22499 0 diode
R22500 N22499 N22500 10
D22500 N22500 0 diode
R22501 N22500 N22501 10
D22501 N22501 0 diode
R22502 N22501 N22502 10
D22502 N22502 0 diode
R22503 N22502 N22503 10
D22503 N22503 0 diode
R22504 N22503 N22504 10
D22504 N22504 0 diode
R22505 N22504 N22505 10
D22505 N22505 0 diode
R22506 N22505 N22506 10
D22506 N22506 0 diode
R22507 N22506 N22507 10
D22507 N22507 0 diode
R22508 N22507 N22508 10
D22508 N22508 0 diode
R22509 N22508 N22509 10
D22509 N22509 0 diode
R22510 N22509 N22510 10
D22510 N22510 0 diode
R22511 N22510 N22511 10
D22511 N22511 0 diode
R22512 N22511 N22512 10
D22512 N22512 0 diode
R22513 N22512 N22513 10
D22513 N22513 0 diode
R22514 N22513 N22514 10
D22514 N22514 0 diode
R22515 N22514 N22515 10
D22515 N22515 0 diode
R22516 N22515 N22516 10
D22516 N22516 0 diode
R22517 N22516 N22517 10
D22517 N22517 0 diode
R22518 N22517 N22518 10
D22518 N22518 0 diode
R22519 N22518 N22519 10
D22519 N22519 0 diode
R22520 N22519 N22520 10
D22520 N22520 0 diode
R22521 N22520 N22521 10
D22521 N22521 0 diode
R22522 N22521 N22522 10
D22522 N22522 0 diode
R22523 N22522 N22523 10
D22523 N22523 0 diode
R22524 N22523 N22524 10
D22524 N22524 0 diode
R22525 N22524 N22525 10
D22525 N22525 0 diode
R22526 N22525 N22526 10
D22526 N22526 0 diode
R22527 N22526 N22527 10
D22527 N22527 0 diode
R22528 N22527 N22528 10
D22528 N22528 0 diode
R22529 N22528 N22529 10
D22529 N22529 0 diode
R22530 N22529 N22530 10
D22530 N22530 0 diode
R22531 N22530 N22531 10
D22531 N22531 0 diode
R22532 N22531 N22532 10
D22532 N22532 0 diode
R22533 N22532 N22533 10
D22533 N22533 0 diode
R22534 N22533 N22534 10
D22534 N22534 0 diode
R22535 N22534 N22535 10
D22535 N22535 0 diode
R22536 N22535 N22536 10
D22536 N22536 0 diode
R22537 N22536 N22537 10
D22537 N22537 0 diode
R22538 N22537 N22538 10
D22538 N22538 0 diode
R22539 N22538 N22539 10
D22539 N22539 0 diode
R22540 N22539 N22540 10
D22540 N22540 0 diode
R22541 N22540 N22541 10
D22541 N22541 0 diode
R22542 N22541 N22542 10
D22542 N22542 0 diode
R22543 N22542 N22543 10
D22543 N22543 0 diode
R22544 N22543 N22544 10
D22544 N22544 0 diode
R22545 N22544 N22545 10
D22545 N22545 0 diode
R22546 N22545 N22546 10
D22546 N22546 0 diode
R22547 N22546 N22547 10
D22547 N22547 0 diode
R22548 N22547 N22548 10
D22548 N22548 0 diode
R22549 N22548 N22549 10
D22549 N22549 0 diode
R22550 N22549 N22550 10
D22550 N22550 0 diode
R22551 N22550 N22551 10
D22551 N22551 0 diode
R22552 N22551 N22552 10
D22552 N22552 0 diode
R22553 N22552 N22553 10
D22553 N22553 0 diode
R22554 N22553 N22554 10
D22554 N22554 0 diode
R22555 N22554 N22555 10
D22555 N22555 0 diode
R22556 N22555 N22556 10
D22556 N22556 0 diode
R22557 N22556 N22557 10
D22557 N22557 0 diode
R22558 N22557 N22558 10
D22558 N22558 0 diode
R22559 N22558 N22559 10
D22559 N22559 0 diode
R22560 N22559 N22560 10
D22560 N22560 0 diode
R22561 N22560 N22561 10
D22561 N22561 0 diode
R22562 N22561 N22562 10
D22562 N22562 0 diode
R22563 N22562 N22563 10
D22563 N22563 0 diode
R22564 N22563 N22564 10
D22564 N22564 0 diode
R22565 N22564 N22565 10
D22565 N22565 0 diode
R22566 N22565 N22566 10
D22566 N22566 0 diode
R22567 N22566 N22567 10
D22567 N22567 0 diode
R22568 N22567 N22568 10
D22568 N22568 0 diode
R22569 N22568 N22569 10
D22569 N22569 0 diode
R22570 N22569 N22570 10
D22570 N22570 0 diode
R22571 N22570 N22571 10
D22571 N22571 0 diode
R22572 N22571 N22572 10
D22572 N22572 0 diode
R22573 N22572 N22573 10
D22573 N22573 0 diode
R22574 N22573 N22574 10
D22574 N22574 0 diode
R22575 N22574 N22575 10
D22575 N22575 0 diode
R22576 N22575 N22576 10
D22576 N22576 0 diode
R22577 N22576 N22577 10
D22577 N22577 0 diode
R22578 N22577 N22578 10
D22578 N22578 0 diode
R22579 N22578 N22579 10
D22579 N22579 0 diode
R22580 N22579 N22580 10
D22580 N22580 0 diode
R22581 N22580 N22581 10
D22581 N22581 0 diode
R22582 N22581 N22582 10
D22582 N22582 0 diode
R22583 N22582 N22583 10
D22583 N22583 0 diode
R22584 N22583 N22584 10
D22584 N22584 0 diode
R22585 N22584 N22585 10
D22585 N22585 0 diode
R22586 N22585 N22586 10
D22586 N22586 0 diode
R22587 N22586 N22587 10
D22587 N22587 0 diode
R22588 N22587 N22588 10
D22588 N22588 0 diode
R22589 N22588 N22589 10
D22589 N22589 0 diode
R22590 N22589 N22590 10
D22590 N22590 0 diode
R22591 N22590 N22591 10
D22591 N22591 0 diode
R22592 N22591 N22592 10
D22592 N22592 0 diode
R22593 N22592 N22593 10
D22593 N22593 0 diode
R22594 N22593 N22594 10
D22594 N22594 0 diode
R22595 N22594 N22595 10
D22595 N22595 0 diode
R22596 N22595 N22596 10
D22596 N22596 0 diode
R22597 N22596 N22597 10
D22597 N22597 0 diode
R22598 N22597 N22598 10
D22598 N22598 0 diode
R22599 N22598 N22599 10
D22599 N22599 0 diode
R22600 N22599 N22600 10
D22600 N22600 0 diode
R22601 N22600 N22601 10
D22601 N22601 0 diode
R22602 N22601 N22602 10
D22602 N22602 0 diode
R22603 N22602 N22603 10
D22603 N22603 0 diode
R22604 N22603 N22604 10
D22604 N22604 0 diode
R22605 N22604 N22605 10
D22605 N22605 0 diode
R22606 N22605 N22606 10
D22606 N22606 0 diode
R22607 N22606 N22607 10
D22607 N22607 0 diode
R22608 N22607 N22608 10
D22608 N22608 0 diode
R22609 N22608 N22609 10
D22609 N22609 0 diode
R22610 N22609 N22610 10
D22610 N22610 0 diode
R22611 N22610 N22611 10
D22611 N22611 0 diode
R22612 N22611 N22612 10
D22612 N22612 0 diode
R22613 N22612 N22613 10
D22613 N22613 0 diode
R22614 N22613 N22614 10
D22614 N22614 0 diode
R22615 N22614 N22615 10
D22615 N22615 0 diode
R22616 N22615 N22616 10
D22616 N22616 0 diode
R22617 N22616 N22617 10
D22617 N22617 0 diode
R22618 N22617 N22618 10
D22618 N22618 0 diode
R22619 N22618 N22619 10
D22619 N22619 0 diode
R22620 N22619 N22620 10
D22620 N22620 0 diode
R22621 N22620 N22621 10
D22621 N22621 0 diode
R22622 N22621 N22622 10
D22622 N22622 0 diode
R22623 N22622 N22623 10
D22623 N22623 0 diode
R22624 N22623 N22624 10
D22624 N22624 0 diode
R22625 N22624 N22625 10
D22625 N22625 0 diode
R22626 N22625 N22626 10
D22626 N22626 0 diode
R22627 N22626 N22627 10
D22627 N22627 0 diode
R22628 N22627 N22628 10
D22628 N22628 0 diode
R22629 N22628 N22629 10
D22629 N22629 0 diode
R22630 N22629 N22630 10
D22630 N22630 0 diode
R22631 N22630 N22631 10
D22631 N22631 0 diode
R22632 N22631 N22632 10
D22632 N22632 0 diode
R22633 N22632 N22633 10
D22633 N22633 0 diode
R22634 N22633 N22634 10
D22634 N22634 0 diode
R22635 N22634 N22635 10
D22635 N22635 0 diode
R22636 N22635 N22636 10
D22636 N22636 0 diode
R22637 N22636 N22637 10
D22637 N22637 0 diode
R22638 N22637 N22638 10
D22638 N22638 0 diode
R22639 N22638 N22639 10
D22639 N22639 0 diode
R22640 N22639 N22640 10
D22640 N22640 0 diode
R22641 N22640 N22641 10
D22641 N22641 0 diode
R22642 N22641 N22642 10
D22642 N22642 0 diode
R22643 N22642 N22643 10
D22643 N22643 0 diode
R22644 N22643 N22644 10
D22644 N22644 0 diode
R22645 N22644 N22645 10
D22645 N22645 0 diode
R22646 N22645 N22646 10
D22646 N22646 0 diode
R22647 N22646 N22647 10
D22647 N22647 0 diode
R22648 N22647 N22648 10
D22648 N22648 0 diode
R22649 N22648 N22649 10
D22649 N22649 0 diode
R22650 N22649 N22650 10
D22650 N22650 0 diode
R22651 N22650 N22651 10
D22651 N22651 0 diode
R22652 N22651 N22652 10
D22652 N22652 0 diode
R22653 N22652 N22653 10
D22653 N22653 0 diode
R22654 N22653 N22654 10
D22654 N22654 0 diode
R22655 N22654 N22655 10
D22655 N22655 0 diode
R22656 N22655 N22656 10
D22656 N22656 0 diode
R22657 N22656 N22657 10
D22657 N22657 0 diode
R22658 N22657 N22658 10
D22658 N22658 0 diode
R22659 N22658 N22659 10
D22659 N22659 0 diode
R22660 N22659 N22660 10
D22660 N22660 0 diode
R22661 N22660 N22661 10
D22661 N22661 0 diode
R22662 N22661 N22662 10
D22662 N22662 0 diode
R22663 N22662 N22663 10
D22663 N22663 0 diode
R22664 N22663 N22664 10
D22664 N22664 0 diode
R22665 N22664 N22665 10
D22665 N22665 0 diode
R22666 N22665 N22666 10
D22666 N22666 0 diode
R22667 N22666 N22667 10
D22667 N22667 0 diode
R22668 N22667 N22668 10
D22668 N22668 0 diode
R22669 N22668 N22669 10
D22669 N22669 0 diode
R22670 N22669 N22670 10
D22670 N22670 0 diode
R22671 N22670 N22671 10
D22671 N22671 0 diode
R22672 N22671 N22672 10
D22672 N22672 0 diode
R22673 N22672 N22673 10
D22673 N22673 0 diode
R22674 N22673 N22674 10
D22674 N22674 0 diode
R22675 N22674 N22675 10
D22675 N22675 0 diode
R22676 N22675 N22676 10
D22676 N22676 0 diode
R22677 N22676 N22677 10
D22677 N22677 0 diode
R22678 N22677 N22678 10
D22678 N22678 0 diode
R22679 N22678 N22679 10
D22679 N22679 0 diode
R22680 N22679 N22680 10
D22680 N22680 0 diode
R22681 N22680 N22681 10
D22681 N22681 0 diode
R22682 N22681 N22682 10
D22682 N22682 0 diode
R22683 N22682 N22683 10
D22683 N22683 0 diode
R22684 N22683 N22684 10
D22684 N22684 0 diode
R22685 N22684 N22685 10
D22685 N22685 0 diode
R22686 N22685 N22686 10
D22686 N22686 0 diode
R22687 N22686 N22687 10
D22687 N22687 0 diode
R22688 N22687 N22688 10
D22688 N22688 0 diode
R22689 N22688 N22689 10
D22689 N22689 0 diode
R22690 N22689 N22690 10
D22690 N22690 0 diode
R22691 N22690 N22691 10
D22691 N22691 0 diode
R22692 N22691 N22692 10
D22692 N22692 0 diode
R22693 N22692 N22693 10
D22693 N22693 0 diode
R22694 N22693 N22694 10
D22694 N22694 0 diode
R22695 N22694 N22695 10
D22695 N22695 0 diode
R22696 N22695 N22696 10
D22696 N22696 0 diode
R22697 N22696 N22697 10
D22697 N22697 0 diode
R22698 N22697 N22698 10
D22698 N22698 0 diode
R22699 N22698 N22699 10
D22699 N22699 0 diode
R22700 N22699 N22700 10
D22700 N22700 0 diode
R22701 N22700 N22701 10
D22701 N22701 0 diode
R22702 N22701 N22702 10
D22702 N22702 0 diode
R22703 N22702 N22703 10
D22703 N22703 0 diode
R22704 N22703 N22704 10
D22704 N22704 0 diode
R22705 N22704 N22705 10
D22705 N22705 0 diode
R22706 N22705 N22706 10
D22706 N22706 0 diode
R22707 N22706 N22707 10
D22707 N22707 0 diode
R22708 N22707 N22708 10
D22708 N22708 0 diode
R22709 N22708 N22709 10
D22709 N22709 0 diode
R22710 N22709 N22710 10
D22710 N22710 0 diode
R22711 N22710 N22711 10
D22711 N22711 0 diode
R22712 N22711 N22712 10
D22712 N22712 0 diode
R22713 N22712 N22713 10
D22713 N22713 0 diode
R22714 N22713 N22714 10
D22714 N22714 0 diode
R22715 N22714 N22715 10
D22715 N22715 0 diode
R22716 N22715 N22716 10
D22716 N22716 0 diode
R22717 N22716 N22717 10
D22717 N22717 0 diode
R22718 N22717 N22718 10
D22718 N22718 0 diode
R22719 N22718 N22719 10
D22719 N22719 0 diode
R22720 N22719 N22720 10
D22720 N22720 0 diode
R22721 N22720 N22721 10
D22721 N22721 0 diode
R22722 N22721 N22722 10
D22722 N22722 0 diode
R22723 N22722 N22723 10
D22723 N22723 0 diode
R22724 N22723 N22724 10
D22724 N22724 0 diode
R22725 N22724 N22725 10
D22725 N22725 0 diode
R22726 N22725 N22726 10
D22726 N22726 0 diode
R22727 N22726 N22727 10
D22727 N22727 0 diode
R22728 N22727 N22728 10
D22728 N22728 0 diode
R22729 N22728 N22729 10
D22729 N22729 0 diode
R22730 N22729 N22730 10
D22730 N22730 0 diode
R22731 N22730 N22731 10
D22731 N22731 0 diode
R22732 N22731 N22732 10
D22732 N22732 0 diode
R22733 N22732 N22733 10
D22733 N22733 0 diode
R22734 N22733 N22734 10
D22734 N22734 0 diode
R22735 N22734 N22735 10
D22735 N22735 0 diode
R22736 N22735 N22736 10
D22736 N22736 0 diode
R22737 N22736 N22737 10
D22737 N22737 0 diode
R22738 N22737 N22738 10
D22738 N22738 0 diode
R22739 N22738 N22739 10
D22739 N22739 0 diode
R22740 N22739 N22740 10
D22740 N22740 0 diode
R22741 N22740 N22741 10
D22741 N22741 0 diode
R22742 N22741 N22742 10
D22742 N22742 0 diode
R22743 N22742 N22743 10
D22743 N22743 0 diode
R22744 N22743 N22744 10
D22744 N22744 0 diode
R22745 N22744 N22745 10
D22745 N22745 0 diode
R22746 N22745 N22746 10
D22746 N22746 0 diode
R22747 N22746 N22747 10
D22747 N22747 0 diode
R22748 N22747 N22748 10
D22748 N22748 0 diode
R22749 N22748 N22749 10
D22749 N22749 0 diode
R22750 N22749 N22750 10
D22750 N22750 0 diode
R22751 N22750 N22751 10
D22751 N22751 0 diode
R22752 N22751 N22752 10
D22752 N22752 0 diode
R22753 N22752 N22753 10
D22753 N22753 0 diode
R22754 N22753 N22754 10
D22754 N22754 0 diode
R22755 N22754 N22755 10
D22755 N22755 0 diode
R22756 N22755 N22756 10
D22756 N22756 0 diode
R22757 N22756 N22757 10
D22757 N22757 0 diode
R22758 N22757 N22758 10
D22758 N22758 0 diode
R22759 N22758 N22759 10
D22759 N22759 0 diode
R22760 N22759 N22760 10
D22760 N22760 0 diode
R22761 N22760 N22761 10
D22761 N22761 0 diode
R22762 N22761 N22762 10
D22762 N22762 0 diode
R22763 N22762 N22763 10
D22763 N22763 0 diode
R22764 N22763 N22764 10
D22764 N22764 0 diode
R22765 N22764 N22765 10
D22765 N22765 0 diode
R22766 N22765 N22766 10
D22766 N22766 0 diode
R22767 N22766 N22767 10
D22767 N22767 0 diode
R22768 N22767 N22768 10
D22768 N22768 0 diode
R22769 N22768 N22769 10
D22769 N22769 0 diode
R22770 N22769 N22770 10
D22770 N22770 0 diode
R22771 N22770 N22771 10
D22771 N22771 0 diode
R22772 N22771 N22772 10
D22772 N22772 0 diode
R22773 N22772 N22773 10
D22773 N22773 0 diode
R22774 N22773 N22774 10
D22774 N22774 0 diode
R22775 N22774 N22775 10
D22775 N22775 0 diode
R22776 N22775 N22776 10
D22776 N22776 0 diode
R22777 N22776 N22777 10
D22777 N22777 0 diode
R22778 N22777 N22778 10
D22778 N22778 0 diode
R22779 N22778 N22779 10
D22779 N22779 0 diode
R22780 N22779 N22780 10
D22780 N22780 0 diode
R22781 N22780 N22781 10
D22781 N22781 0 diode
R22782 N22781 N22782 10
D22782 N22782 0 diode
R22783 N22782 N22783 10
D22783 N22783 0 diode
R22784 N22783 N22784 10
D22784 N22784 0 diode
R22785 N22784 N22785 10
D22785 N22785 0 diode
R22786 N22785 N22786 10
D22786 N22786 0 diode
R22787 N22786 N22787 10
D22787 N22787 0 diode
R22788 N22787 N22788 10
D22788 N22788 0 diode
R22789 N22788 N22789 10
D22789 N22789 0 diode
R22790 N22789 N22790 10
D22790 N22790 0 diode
R22791 N22790 N22791 10
D22791 N22791 0 diode
R22792 N22791 N22792 10
D22792 N22792 0 diode
R22793 N22792 N22793 10
D22793 N22793 0 diode
R22794 N22793 N22794 10
D22794 N22794 0 diode
R22795 N22794 N22795 10
D22795 N22795 0 diode
R22796 N22795 N22796 10
D22796 N22796 0 diode
R22797 N22796 N22797 10
D22797 N22797 0 diode
R22798 N22797 N22798 10
D22798 N22798 0 diode
R22799 N22798 N22799 10
D22799 N22799 0 diode
R22800 N22799 N22800 10
D22800 N22800 0 diode
R22801 N22800 N22801 10
D22801 N22801 0 diode
R22802 N22801 N22802 10
D22802 N22802 0 diode
R22803 N22802 N22803 10
D22803 N22803 0 diode
R22804 N22803 N22804 10
D22804 N22804 0 diode
R22805 N22804 N22805 10
D22805 N22805 0 diode
R22806 N22805 N22806 10
D22806 N22806 0 diode
R22807 N22806 N22807 10
D22807 N22807 0 diode
R22808 N22807 N22808 10
D22808 N22808 0 diode
R22809 N22808 N22809 10
D22809 N22809 0 diode
R22810 N22809 N22810 10
D22810 N22810 0 diode
R22811 N22810 N22811 10
D22811 N22811 0 diode
R22812 N22811 N22812 10
D22812 N22812 0 diode
R22813 N22812 N22813 10
D22813 N22813 0 diode
R22814 N22813 N22814 10
D22814 N22814 0 diode
R22815 N22814 N22815 10
D22815 N22815 0 diode
R22816 N22815 N22816 10
D22816 N22816 0 diode
R22817 N22816 N22817 10
D22817 N22817 0 diode
R22818 N22817 N22818 10
D22818 N22818 0 diode
R22819 N22818 N22819 10
D22819 N22819 0 diode
R22820 N22819 N22820 10
D22820 N22820 0 diode
R22821 N22820 N22821 10
D22821 N22821 0 diode
R22822 N22821 N22822 10
D22822 N22822 0 diode
R22823 N22822 N22823 10
D22823 N22823 0 diode
R22824 N22823 N22824 10
D22824 N22824 0 diode
R22825 N22824 N22825 10
D22825 N22825 0 diode
R22826 N22825 N22826 10
D22826 N22826 0 diode
R22827 N22826 N22827 10
D22827 N22827 0 diode
R22828 N22827 N22828 10
D22828 N22828 0 diode
R22829 N22828 N22829 10
D22829 N22829 0 diode
R22830 N22829 N22830 10
D22830 N22830 0 diode
R22831 N22830 N22831 10
D22831 N22831 0 diode
R22832 N22831 N22832 10
D22832 N22832 0 diode
R22833 N22832 N22833 10
D22833 N22833 0 diode
R22834 N22833 N22834 10
D22834 N22834 0 diode
R22835 N22834 N22835 10
D22835 N22835 0 diode
R22836 N22835 N22836 10
D22836 N22836 0 diode
R22837 N22836 N22837 10
D22837 N22837 0 diode
R22838 N22837 N22838 10
D22838 N22838 0 diode
R22839 N22838 N22839 10
D22839 N22839 0 diode
R22840 N22839 N22840 10
D22840 N22840 0 diode
R22841 N22840 N22841 10
D22841 N22841 0 diode
R22842 N22841 N22842 10
D22842 N22842 0 diode
R22843 N22842 N22843 10
D22843 N22843 0 diode
R22844 N22843 N22844 10
D22844 N22844 0 diode
R22845 N22844 N22845 10
D22845 N22845 0 diode
R22846 N22845 N22846 10
D22846 N22846 0 diode
R22847 N22846 N22847 10
D22847 N22847 0 diode
R22848 N22847 N22848 10
D22848 N22848 0 diode
R22849 N22848 N22849 10
D22849 N22849 0 diode
R22850 N22849 N22850 10
D22850 N22850 0 diode
R22851 N22850 N22851 10
D22851 N22851 0 diode
R22852 N22851 N22852 10
D22852 N22852 0 diode
R22853 N22852 N22853 10
D22853 N22853 0 diode
R22854 N22853 N22854 10
D22854 N22854 0 diode
R22855 N22854 N22855 10
D22855 N22855 0 diode
R22856 N22855 N22856 10
D22856 N22856 0 diode
R22857 N22856 N22857 10
D22857 N22857 0 diode
R22858 N22857 N22858 10
D22858 N22858 0 diode
R22859 N22858 N22859 10
D22859 N22859 0 diode
R22860 N22859 N22860 10
D22860 N22860 0 diode
R22861 N22860 N22861 10
D22861 N22861 0 diode
R22862 N22861 N22862 10
D22862 N22862 0 diode
R22863 N22862 N22863 10
D22863 N22863 0 diode
R22864 N22863 N22864 10
D22864 N22864 0 diode
R22865 N22864 N22865 10
D22865 N22865 0 diode
R22866 N22865 N22866 10
D22866 N22866 0 diode
R22867 N22866 N22867 10
D22867 N22867 0 diode
R22868 N22867 N22868 10
D22868 N22868 0 diode
R22869 N22868 N22869 10
D22869 N22869 0 diode
R22870 N22869 N22870 10
D22870 N22870 0 diode
R22871 N22870 N22871 10
D22871 N22871 0 diode
R22872 N22871 N22872 10
D22872 N22872 0 diode
R22873 N22872 N22873 10
D22873 N22873 0 diode
R22874 N22873 N22874 10
D22874 N22874 0 diode
R22875 N22874 N22875 10
D22875 N22875 0 diode
R22876 N22875 N22876 10
D22876 N22876 0 diode
R22877 N22876 N22877 10
D22877 N22877 0 diode
R22878 N22877 N22878 10
D22878 N22878 0 diode
R22879 N22878 N22879 10
D22879 N22879 0 diode
R22880 N22879 N22880 10
D22880 N22880 0 diode
R22881 N22880 N22881 10
D22881 N22881 0 diode
R22882 N22881 N22882 10
D22882 N22882 0 diode
R22883 N22882 N22883 10
D22883 N22883 0 diode
R22884 N22883 N22884 10
D22884 N22884 0 diode
R22885 N22884 N22885 10
D22885 N22885 0 diode
R22886 N22885 N22886 10
D22886 N22886 0 diode
R22887 N22886 N22887 10
D22887 N22887 0 diode
R22888 N22887 N22888 10
D22888 N22888 0 diode
R22889 N22888 N22889 10
D22889 N22889 0 diode
R22890 N22889 N22890 10
D22890 N22890 0 diode
R22891 N22890 N22891 10
D22891 N22891 0 diode
R22892 N22891 N22892 10
D22892 N22892 0 diode
R22893 N22892 N22893 10
D22893 N22893 0 diode
R22894 N22893 N22894 10
D22894 N22894 0 diode
R22895 N22894 N22895 10
D22895 N22895 0 diode
R22896 N22895 N22896 10
D22896 N22896 0 diode
R22897 N22896 N22897 10
D22897 N22897 0 diode
R22898 N22897 N22898 10
D22898 N22898 0 diode
R22899 N22898 N22899 10
D22899 N22899 0 diode
R22900 N22899 N22900 10
D22900 N22900 0 diode
R22901 N22900 N22901 10
D22901 N22901 0 diode
R22902 N22901 N22902 10
D22902 N22902 0 diode
R22903 N22902 N22903 10
D22903 N22903 0 diode
R22904 N22903 N22904 10
D22904 N22904 0 diode
R22905 N22904 N22905 10
D22905 N22905 0 diode
R22906 N22905 N22906 10
D22906 N22906 0 diode
R22907 N22906 N22907 10
D22907 N22907 0 diode
R22908 N22907 N22908 10
D22908 N22908 0 diode
R22909 N22908 N22909 10
D22909 N22909 0 diode
R22910 N22909 N22910 10
D22910 N22910 0 diode
R22911 N22910 N22911 10
D22911 N22911 0 diode
R22912 N22911 N22912 10
D22912 N22912 0 diode
R22913 N22912 N22913 10
D22913 N22913 0 diode
R22914 N22913 N22914 10
D22914 N22914 0 diode
R22915 N22914 N22915 10
D22915 N22915 0 diode
R22916 N22915 N22916 10
D22916 N22916 0 diode
R22917 N22916 N22917 10
D22917 N22917 0 diode
R22918 N22917 N22918 10
D22918 N22918 0 diode
R22919 N22918 N22919 10
D22919 N22919 0 diode
R22920 N22919 N22920 10
D22920 N22920 0 diode
R22921 N22920 N22921 10
D22921 N22921 0 diode
R22922 N22921 N22922 10
D22922 N22922 0 diode
R22923 N22922 N22923 10
D22923 N22923 0 diode
R22924 N22923 N22924 10
D22924 N22924 0 diode
R22925 N22924 N22925 10
D22925 N22925 0 diode
R22926 N22925 N22926 10
D22926 N22926 0 diode
R22927 N22926 N22927 10
D22927 N22927 0 diode
R22928 N22927 N22928 10
D22928 N22928 0 diode
R22929 N22928 N22929 10
D22929 N22929 0 diode
R22930 N22929 N22930 10
D22930 N22930 0 diode
R22931 N22930 N22931 10
D22931 N22931 0 diode
R22932 N22931 N22932 10
D22932 N22932 0 diode
R22933 N22932 N22933 10
D22933 N22933 0 diode
R22934 N22933 N22934 10
D22934 N22934 0 diode
R22935 N22934 N22935 10
D22935 N22935 0 diode
R22936 N22935 N22936 10
D22936 N22936 0 diode
R22937 N22936 N22937 10
D22937 N22937 0 diode
R22938 N22937 N22938 10
D22938 N22938 0 diode
R22939 N22938 N22939 10
D22939 N22939 0 diode
R22940 N22939 N22940 10
D22940 N22940 0 diode
R22941 N22940 N22941 10
D22941 N22941 0 diode
R22942 N22941 N22942 10
D22942 N22942 0 diode
R22943 N22942 N22943 10
D22943 N22943 0 diode
R22944 N22943 N22944 10
D22944 N22944 0 diode
R22945 N22944 N22945 10
D22945 N22945 0 diode
R22946 N22945 N22946 10
D22946 N22946 0 diode
R22947 N22946 N22947 10
D22947 N22947 0 diode
R22948 N22947 N22948 10
D22948 N22948 0 diode
R22949 N22948 N22949 10
D22949 N22949 0 diode
R22950 N22949 N22950 10
D22950 N22950 0 diode
R22951 N22950 N22951 10
D22951 N22951 0 diode
R22952 N22951 N22952 10
D22952 N22952 0 diode
R22953 N22952 N22953 10
D22953 N22953 0 diode
R22954 N22953 N22954 10
D22954 N22954 0 diode
R22955 N22954 N22955 10
D22955 N22955 0 diode
R22956 N22955 N22956 10
D22956 N22956 0 diode
R22957 N22956 N22957 10
D22957 N22957 0 diode
R22958 N22957 N22958 10
D22958 N22958 0 diode
R22959 N22958 N22959 10
D22959 N22959 0 diode
R22960 N22959 N22960 10
D22960 N22960 0 diode
R22961 N22960 N22961 10
D22961 N22961 0 diode
R22962 N22961 N22962 10
D22962 N22962 0 diode
R22963 N22962 N22963 10
D22963 N22963 0 diode
R22964 N22963 N22964 10
D22964 N22964 0 diode
R22965 N22964 N22965 10
D22965 N22965 0 diode
R22966 N22965 N22966 10
D22966 N22966 0 diode
R22967 N22966 N22967 10
D22967 N22967 0 diode
R22968 N22967 N22968 10
D22968 N22968 0 diode
R22969 N22968 N22969 10
D22969 N22969 0 diode
R22970 N22969 N22970 10
D22970 N22970 0 diode
R22971 N22970 N22971 10
D22971 N22971 0 diode
R22972 N22971 N22972 10
D22972 N22972 0 diode
R22973 N22972 N22973 10
D22973 N22973 0 diode
R22974 N22973 N22974 10
D22974 N22974 0 diode
R22975 N22974 N22975 10
D22975 N22975 0 diode
R22976 N22975 N22976 10
D22976 N22976 0 diode
R22977 N22976 N22977 10
D22977 N22977 0 diode
R22978 N22977 N22978 10
D22978 N22978 0 diode
R22979 N22978 N22979 10
D22979 N22979 0 diode
R22980 N22979 N22980 10
D22980 N22980 0 diode
R22981 N22980 N22981 10
D22981 N22981 0 diode
R22982 N22981 N22982 10
D22982 N22982 0 diode
R22983 N22982 N22983 10
D22983 N22983 0 diode
R22984 N22983 N22984 10
D22984 N22984 0 diode
R22985 N22984 N22985 10
D22985 N22985 0 diode
R22986 N22985 N22986 10
D22986 N22986 0 diode
R22987 N22986 N22987 10
D22987 N22987 0 diode
R22988 N22987 N22988 10
D22988 N22988 0 diode
R22989 N22988 N22989 10
D22989 N22989 0 diode
R22990 N22989 N22990 10
D22990 N22990 0 diode
R22991 N22990 N22991 10
D22991 N22991 0 diode
R22992 N22991 N22992 10
D22992 N22992 0 diode
R22993 N22992 N22993 10
D22993 N22993 0 diode
R22994 N22993 N22994 10
D22994 N22994 0 diode
R22995 N22994 N22995 10
D22995 N22995 0 diode
R22996 N22995 N22996 10
D22996 N22996 0 diode
R22997 N22996 N22997 10
D22997 N22997 0 diode
R22998 N22997 N22998 10
D22998 N22998 0 diode
R22999 N22998 N22999 10
D22999 N22999 0 diode
R23000 N22999 N23000 10
D23000 N23000 0 diode
R23001 N23000 N23001 10
D23001 N23001 0 diode
R23002 N23001 N23002 10
D23002 N23002 0 diode
R23003 N23002 N23003 10
D23003 N23003 0 diode
R23004 N23003 N23004 10
D23004 N23004 0 diode
R23005 N23004 N23005 10
D23005 N23005 0 diode
R23006 N23005 N23006 10
D23006 N23006 0 diode
R23007 N23006 N23007 10
D23007 N23007 0 diode
R23008 N23007 N23008 10
D23008 N23008 0 diode
R23009 N23008 N23009 10
D23009 N23009 0 diode
R23010 N23009 N23010 10
D23010 N23010 0 diode
R23011 N23010 N23011 10
D23011 N23011 0 diode
R23012 N23011 N23012 10
D23012 N23012 0 diode
R23013 N23012 N23013 10
D23013 N23013 0 diode
R23014 N23013 N23014 10
D23014 N23014 0 diode
R23015 N23014 N23015 10
D23015 N23015 0 diode
R23016 N23015 N23016 10
D23016 N23016 0 diode
R23017 N23016 N23017 10
D23017 N23017 0 diode
R23018 N23017 N23018 10
D23018 N23018 0 diode
R23019 N23018 N23019 10
D23019 N23019 0 diode
R23020 N23019 N23020 10
D23020 N23020 0 diode
R23021 N23020 N23021 10
D23021 N23021 0 diode
R23022 N23021 N23022 10
D23022 N23022 0 diode
R23023 N23022 N23023 10
D23023 N23023 0 diode
R23024 N23023 N23024 10
D23024 N23024 0 diode
R23025 N23024 N23025 10
D23025 N23025 0 diode
R23026 N23025 N23026 10
D23026 N23026 0 diode
R23027 N23026 N23027 10
D23027 N23027 0 diode
R23028 N23027 N23028 10
D23028 N23028 0 diode
R23029 N23028 N23029 10
D23029 N23029 0 diode
R23030 N23029 N23030 10
D23030 N23030 0 diode
R23031 N23030 N23031 10
D23031 N23031 0 diode
R23032 N23031 N23032 10
D23032 N23032 0 diode
R23033 N23032 N23033 10
D23033 N23033 0 diode
R23034 N23033 N23034 10
D23034 N23034 0 diode
R23035 N23034 N23035 10
D23035 N23035 0 diode
R23036 N23035 N23036 10
D23036 N23036 0 diode
R23037 N23036 N23037 10
D23037 N23037 0 diode
R23038 N23037 N23038 10
D23038 N23038 0 diode
R23039 N23038 N23039 10
D23039 N23039 0 diode
R23040 N23039 N23040 10
D23040 N23040 0 diode
R23041 N23040 N23041 10
D23041 N23041 0 diode
R23042 N23041 N23042 10
D23042 N23042 0 diode
R23043 N23042 N23043 10
D23043 N23043 0 diode
R23044 N23043 N23044 10
D23044 N23044 0 diode
R23045 N23044 N23045 10
D23045 N23045 0 diode
R23046 N23045 N23046 10
D23046 N23046 0 diode
R23047 N23046 N23047 10
D23047 N23047 0 diode
R23048 N23047 N23048 10
D23048 N23048 0 diode
R23049 N23048 N23049 10
D23049 N23049 0 diode
R23050 N23049 N23050 10
D23050 N23050 0 diode
R23051 N23050 N23051 10
D23051 N23051 0 diode
R23052 N23051 N23052 10
D23052 N23052 0 diode
R23053 N23052 N23053 10
D23053 N23053 0 diode
R23054 N23053 N23054 10
D23054 N23054 0 diode
R23055 N23054 N23055 10
D23055 N23055 0 diode
R23056 N23055 N23056 10
D23056 N23056 0 diode
R23057 N23056 N23057 10
D23057 N23057 0 diode
R23058 N23057 N23058 10
D23058 N23058 0 diode
R23059 N23058 N23059 10
D23059 N23059 0 diode
R23060 N23059 N23060 10
D23060 N23060 0 diode
R23061 N23060 N23061 10
D23061 N23061 0 diode
R23062 N23061 N23062 10
D23062 N23062 0 diode
R23063 N23062 N23063 10
D23063 N23063 0 diode
R23064 N23063 N23064 10
D23064 N23064 0 diode
R23065 N23064 N23065 10
D23065 N23065 0 diode
R23066 N23065 N23066 10
D23066 N23066 0 diode
R23067 N23066 N23067 10
D23067 N23067 0 diode
R23068 N23067 N23068 10
D23068 N23068 0 diode
R23069 N23068 N23069 10
D23069 N23069 0 diode
R23070 N23069 N23070 10
D23070 N23070 0 diode
R23071 N23070 N23071 10
D23071 N23071 0 diode
R23072 N23071 N23072 10
D23072 N23072 0 diode
R23073 N23072 N23073 10
D23073 N23073 0 diode
R23074 N23073 N23074 10
D23074 N23074 0 diode
R23075 N23074 N23075 10
D23075 N23075 0 diode
R23076 N23075 N23076 10
D23076 N23076 0 diode
R23077 N23076 N23077 10
D23077 N23077 0 diode
R23078 N23077 N23078 10
D23078 N23078 0 diode
R23079 N23078 N23079 10
D23079 N23079 0 diode
R23080 N23079 N23080 10
D23080 N23080 0 diode
R23081 N23080 N23081 10
D23081 N23081 0 diode
R23082 N23081 N23082 10
D23082 N23082 0 diode
R23083 N23082 N23083 10
D23083 N23083 0 diode
R23084 N23083 N23084 10
D23084 N23084 0 diode
R23085 N23084 N23085 10
D23085 N23085 0 diode
R23086 N23085 N23086 10
D23086 N23086 0 diode
R23087 N23086 N23087 10
D23087 N23087 0 diode
R23088 N23087 N23088 10
D23088 N23088 0 diode
R23089 N23088 N23089 10
D23089 N23089 0 diode
R23090 N23089 N23090 10
D23090 N23090 0 diode
R23091 N23090 N23091 10
D23091 N23091 0 diode
R23092 N23091 N23092 10
D23092 N23092 0 diode
R23093 N23092 N23093 10
D23093 N23093 0 diode
R23094 N23093 N23094 10
D23094 N23094 0 diode
R23095 N23094 N23095 10
D23095 N23095 0 diode
R23096 N23095 N23096 10
D23096 N23096 0 diode
R23097 N23096 N23097 10
D23097 N23097 0 diode
R23098 N23097 N23098 10
D23098 N23098 0 diode
R23099 N23098 N23099 10
D23099 N23099 0 diode
R23100 N23099 N23100 10
D23100 N23100 0 diode
R23101 N23100 N23101 10
D23101 N23101 0 diode
R23102 N23101 N23102 10
D23102 N23102 0 diode
R23103 N23102 N23103 10
D23103 N23103 0 diode
R23104 N23103 N23104 10
D23104 N23104 0 diode
R23105 N23104 N23105 10
D23105 N23105 0 diode
R23106 N23105 N23106 10
D23106 N23106 0 diode
R23107 N23106 N23107 10
D23107 N23107 0 diode
R23108 N23107 N23108 10
D23108 N23108 0 diode
R23109 N23108 N23109 10
D23109 N23109 0 diode
R23110 N23109 N23110 10
D23110 N23110 0 diode
R23111 N23110 N23111 10
D23111 N23111 0 diode
R23112 N23111 N23112 10
D23112 N23112 0 diode
R23113 N23112 N23113 10
D23113 N23113 0 diode
R23114 N23113 N23114 10
D23114 N23114 0 diode
R23115 N23114 N23115 10
D23115 N23115 0 diode
R23116 N23115 N23116 10
D23116 N23116 0 diode
R23117 N23116 N23117 10
D23117 N23117 0 diode
R23118 N23117 N23118 10
D23118 N23118 0 diode
R23119 N23118 N23119 10
D23119 N23119 0 diode
R23120 N23119 N23120 10
D23120 N23120 0 diode
R23121 N23120 N23121 10
D23121 N23121 0 diode
R23122 N23121 N23122 10
D23122 N23122 0 diode
R23123 N23122 N23123 10
D23123 N23123 0 diode
R23124 N23123 N23124 10
D23124 N23124 0 diode
R23125 N23124 N23125 10
D23125 N23125 0 diode
R23126 N23125 N23126 10
D23126 N23126 0 diode
R23127 N23126 N23127 10
D23127 N23127 0 diode
R23128 N23127 N23128 10
D23128 N23128 0 diode
R23129 N23128 N23129 10
D23129 N23129 0 diode
R23130 N23129 N23130 10
D23130 N23130 0 diode
R23131 N23130 N23131 10
D23131 N23131 0 diode
R23132 N23131 N23132 10
D23132 N23132 0 diode
R23133 N23132 N23133 10
D23133 N23133 0 diode
R23134 N23133 N23134 10
D23134 N23134 0 diode
R23135 N23134 N23135 10
D23135 N23135 0 diode
R23136 N23135 N23136 10
D23136 N23136 0 diode
R23137 N23136 N23137 10
D23137 N23137 0 diode
R23138 N23137 N23138 10
D23138 N23138 0 diode
R23139 N23138 N23139 10
D23139 N23139 0 diode
R23140 N23139 N23140 10
D23140 N23140 0 diode
R23141 N23140 N23141 10
D23141 N23141 0 diode
R23142 N23141 N23142 10
D23142 N23142 0 diode
R23143 N23142 N23143 10
D23143 N23143 0 diode
R23144 N23143 N23144 10
D23144 N23144 0 diode
R23145 N23144 N23145 10
D23145 N23145 0 diode
R23146 N23145 N23146 10
D23146 N23146 0 diode
R23147 N23146 N23147 10
D23147 N23147 0 diode
R23148 N23147 N23148 10
D23148 N23148 0 diode
R23149 N23148 N23149 10
D23149 N23149 0 diode
R23150 N23149 N23150 10
D23150 N23150 0 diode
R23151 N23150 N23151 10
D23151 N23151 0 diode
R23152 N23151 N23152 10
D23152 N23152 0 diode
R23153 N23152 N23153 10
D23153 N23153 0 diode
R23154 N23153 N23154 10
D23154 N23154 0 diode
R23155 N23154 N23155 10
D23155 N23155 0 diode
R23156 N23155 N23156 10
D23156 N23156 0 diode
R23157 N23156 N23157 10
D23157 N23157 0 diode
R23158 N23157 N23158 10
D23158 N23158 0 diode
R23159 N23158 N23159 10
D23159 N23159 0 diode
R23160 N23159 N23160 10
D23160 N23160 0 diode
R23161 N23160 N23161 10
D23161 N23161 0 diode
R23162 N23161 N23162 10
D23162 N23162 0 diode
R23163 N23162 N23163 10
D23163 N23163 0 diode
R23164 N23163 N23164 10
D23164 N23164 0 diode
R23165 N23164 N23165 10
D23165 N23165 0 diode
R23166 N23165 N23166 10
D23166 N23166 0 diode
R23167 N23166 N23167 10
D23167 N23167 0 diode
R23168 N23167 N23168 10
D23168 N23168 0 diode
R23169 N23168 N23169 10
D23169 N23169 0 diode
R23170 N23169 N23170 10
D23170 N23170 0 diode
R23171 N23170 N23171 10
D23171 N23171 0 diode
R23172 N23171 N23172 10
D23172 N23172 0 diode
R23173 N23172 N23173 10
D23173 N23173 0 diode
R23174 N23173 N23174 10
D23174 N23174 0 diode
R23175 N23174 N23175 10
D23175 N23175 0 diode
R23176 N23175 N23176 10
D23176 N23176 0 diode
R23177 N23176 N23177 10
D23177 N23177 0 diode
R23178 N23177 N23178 10
D23178 N23178 0 diode
R23179 N23178 N23179 10
D23179 N23179 0 diode
R23180 N23179 N23180 10
D23180 N23180 0 diode
R23181 N23180 N23181 10
D23181 N23181 0 diode
R23182 N23181 N23182 10
D23182 N23182 0 diode
R23183 N23182 N23183 10
D23183 N23183 0 diode
R23184 N23183 N23184 10
D23184 N23184 0 diode
R23185 N23184 N23185 10
D23185 N23185 0 diode
R23186 N23185 N23186 10
D23186 N23186 0 diode
R23187 N23186 N23187 10
D23187 N23187 0 diode
R23188 N23187 N23188 10
D23188 N23188 0 diode
R23189 N23188 N23189 10
D23189 N23189 0 diode
R23190 N23189 N23190 10
D23190 N23190 0 diode
R23191 N23190 N23191 10
D23191 N23191 0 diode
R23192 N23191 N23192 10
D23192 N23192 0 diode
R23193 N23192 N23193 10
D23193 N23193 0 diode
R23194 N23193 N23194 10
D23194 N23194 0 diode
R23195 N23194 N23195 10
D23195 N23195 0 diode
R23196 N23195 N23196 10
D23196 N23196 0 diode
R23197 N23196 N23197 10
D23197 N23197 0 diode
R23198 N23197 N23198 10
D23198 N23198 0 diode
R23199 N23198 N23199 10
D23199 N23199 0 diode
R23200 N23199 N23200 10
D23200 N23200 0 diode
R23201 N23200 N23201 10
D23201 N23201 0 diode
R23202 N23201 N23202 10
D23202 N23202 0 diode
R23203 N23202 N23203 10
D23203 N23203 0 diode
R23204 N23203 N23204 10
D23204 N23204 0 diode
R23205 N23204 N23205 10
D23205 N23205 0 diode
R23206 N23205 N23206 10
D23206 N23206 0 diode
R23207 N23206 N23207 10
D23207 N23207 0 diode
R23208 N23207 N23208 10
D23208 N23208 0 diode
R23209 N23208 N23209 10
D23209 N23209 0 diode
R23210 N23209 N23210 10
D23210 N23210 0 diode
R23211 N23210 N23211 10
D23211 N23211 0 diode
R23212 N23211 N23212 10
D23212 N23212 0 diode
R23213 N23212 N23213 10
D23213 N23213 0 diode
R23214 N23213 N23214 10
D23214 N23214 0 diode
R23215 N23214 N23215 10
D23215 N23215 0 diode
R23216 N23215 N23216 10
D23216 N23216 0 diode
R23217 N23216 N23217 10
D23217 N23217 0 diode
R23218 N23217 N23218 10
D23218 N23218 0 diode
R23219 N23218 N23219 10
D23219 N23219 0 diode
R23220 N23219 N23220 10
D23220 N23220 0 diode
R23221 N23220 N23221 10
D23221 N23221 0 diode
R23222 N23221 N23222 10
D23222 N23222 0 diode
R23223 N23222 N23223 10
D23223 N23223 0 diode
R23224 N23223 N23224 10
D23224 N23224 0 diode
R23225 N23224 N23225 10
D23225 N23225 0 diode
R23226 N23225 N23226 10
D23226 N23226 0 diode
R23227 N23226 N23227 10
D23227 N23227 0 diode
R23228 N23227 N23228 10
D23228 N23228 0 diode
R23229 N23228 N23229 10
D23229 N23229 0 diode
R23230 N23229 N23230 10
D23230 N23230 0 diode
R23231 N23230 N23231 10
D23231 N23231 0 diode
R23232 N23231 N23232 10
D23232 N23232 0 diode
R23233 N23232 N23233 10
D23233 N23233 0 diode
R23234 N23233 N23234 10
D23234 N23234 0 diode
R23235 N23234 N23235 10
D23235 N23235 0 diode
R23236 N23235 N23236 10
D23236 N23236 0 diode
R23237 N23236 N23237 10
D23237 N23237 0 diode
R23238 N23237 N23238 10
D23238 N23238 0 diode
R23239 N23238 N23239 10
D23239 N23239 0 diode
R23240 N23239 N23240 10
D23240 N23240 0 diode
R23241 N23240 N23241 10
D23241 N23241 0 diode
R23242 N23241 N23242 10
D23242 N23242 0 diode
R23243 N23242 N23243 10
D23243 N23243 0 diode
R23244 N23243 N23244 10
D23244 N23244 0 diode
R23245 N23244 N23245 10
D23245 N23245 0 diode
R23246 N23245 N23246 10
D23246 N23246 0 diode
R23247 N23246 N23247 10
D23247 N23247 0 diode
R23248 N23247 N23248 10
D23248 N23248 0 diode
R23249 N23248 N23249 10
D23249 N23249 0 diode
R23250 N23249 N23250 10
D23250 N23250 0 diode
R23251 N23250 N23251 10
D23251 N23251 0 diode
R23252 N23251 N23252 10
D23252 N23252 0 diode
R23253 N23252 N23253 10
D23253 N23253 0 diode
R23254 N23253 N23254 10
D23254 N23254 0 diode
R23255 N23254 N23255 10
D23255 N23255 0 diode
R23256 N23255 N23256 10
D23256 N23256 0 diode
R23257 N23256 N23257 10
D23257 N23257 0 diode
R23258 N23257 N23258 10
D23258 N23258 0 diode
R23259 N23258 N23259 10
D23259 N23259 0 diode
R23260 N23259 N23260 10
D23260 N23260 0 diode
R23261 N23260 N23261 10
D23261 N23261 0 diode
R23262 N23261 N23262 10
D23262 N23262 0 diode
R23263 N23262 N23263 10
D23263 N23263 0 diode
R23264 N23263 N23264 10
D23264 N23264 0 diode
R23265 N23264 N23265 10
D23265 N23265 0 diode
R23266 N23265 N23266 10
D23266 N23266 0 diode
R23267 N23266 N23267 10
D23267 N23267 0 diode
R23268 N23267 N23268 10
D23268 N23268 0 diode
R23269 N23268 N23269 10
D23269 N23269 0 diode
R23270 N23269 N23270 10
D23270 N23270 0 diode
R23271 N23270 N23271 10
D23271 N23271 0 diode
R23272 N23271 N23272 10
D23272 N23272 0 diode
R23273 N23272 N23273 10
D23273 N23273 0 diode
R23274 N23273 N23274 10
D23274 N23274 0 diode
R23275 N23274 N23275 10
D23275 N23275 0 diode
R23276 N23275 N23276 10
D23276 N23276 0 diode
R23277 N23276 N23277 10
D23277 N23277 0 diode
R23278 N23277 N23278 10
D23278 N23278 0 diode
R23279 N23278 N23279 10
D23279 N23279 0 diode
R23280 N23279 N23280 10
D23280 N23280 0 diode
R23281 N23280 N23281 10
D23281 N23281 0 diode
R23282 N23281 N23282 10
D23282 N23282 0 diode
R23283 N23282 N23283 10
D23283 N23283 0 diode
R23284 N23283 N23284 10
D23284 N23284 0 diode
R23285 N23284 N23285 10
D23285 N23285 0 diode
R23286 N23285 N23286 10
D23286 N23286 0 diode
R23287 N23286 N23287 10
D23287 N23287 0 diode
R23288 N23287 N23288 10
D23288 N23288 0 diode
R23289 N23288 N23289 10
D23289 N23289 0 diode
R23290 N23289 N23290 10
D23290 N23290 0 diode
R23291 N23290 N23291 10
D23291 N23291 0 diode
R23292 N23291 N23292 10
D23292 N23292 0 diode
R23293 N23292 N23293 10
D23293 N23293 0 diode
R23294 N23293 N23294 10
D23294 N23294 0 diode
R23295 N23294 N23295 10
D23295 N23295 0 diode
R23296 N23295 N23296 10
D23296 N23296 0 diode
R23297 N23296 N23297 10
D23297 N23297 0 diode
R23298 N23297 N23298 10
D23298 N23298 0 diode
R23299 N23298 N23299 10
D23299 N23299 0 diode
R23300 N23299 N23300 10
D23300 N23300 0 diode
R23301 N23300 N23301 10
D23301 N23301 0 diode
R23302 N23301 N23302 10
D23302 N23302 0 diode
R23303 N23302 N23303 10
D23303 N23303 0 diode
R23304 N23303 N23304 10
D23304 N23304 0 diode
R23305 N23304 N23305 10
D23305 N23305 0 diode
R23306 N23305 N23306 10
D23306 N23306 0 diode
R23307 N23306 N23307 10
D23307 N23307 0 diode
R23308 N23307 N23308 10
D23308 N23308 0 diode
R23309 N23308 N23309 10
D23309 N23309 0 diode
R23310 N23309 N23310 10
D23310 N23310 0 diode
R23311 N23310 N23311 10
D23311 N23311 0 diode
R23312 N23311 N23312 10
D23312 N23312 0 diode
R23313 N23312 N23313 10
D23313 N23313 0 diode
R23314 N23313 N23314 10
D23314 N23314 0 diode
R23315 N23314 N23315 10
D23315 N23315 0 diode
R23316 N23315 N23316 10
D23316 N23316 0 diode
R23317 N23316 N23317 10
D23317 N23317 0 diode
R23318 N23317 N23318 10
D23318 N23318 0 diode
R23319 N23318 N23319 10
D23319 N23319 0 diode
R23320 N23319 N23320 10
D23320 N23320 0 diode
R23321 N23320 N23321 10
D23321 N23321 0 diode
R23322 N23321 N23322 10
D23322 N23322 0 diode
R23323 N23322 N23323 10
D23323 N23323 0 diode
R23324 N23323 N23324 10
D23324 N23324 0 diode
R23325 N23324 N23325 10
D23325 N23325 0 diode
R23326 N23325 N23326 10
D23326 N23326 0 diode
R23327 N23326 N23327 10
D23327 N23327 0 diode
R23328 N23327 N23328 10
D23328 N23328 0 diode
R23329 N23328 N23329 10
D23329 N23329 0 diode
R23330 N23329 N23330 10
D23330 N23330 0 diode
R23331 N23330 N23331 10
D23331 N23331 0 diode
R23332 N23331 N23332 10
D23332 N23332 0 diode
R23333 N23332 N23333 10
D23333 N23333 0 diode
R23334 N23333 N23334 10
D23334 N23334 0 diode
R23335 N23334 N23335 10
D23335 N23335 0 diode
R23336 N23335 N23336 10
D23336 N23336 0 diode
R23337 N23336 N23337 10
D23337 N23337 0 diode
R23338 N23337 N23338 10
D23338 N23338 0 diode
R23339 N23338 N23339 10
D23339 N23339 0 diode
R23340 N23339 N23340 10
D23340 N23340 0 diode
R23341 N23340 N23341 10
D23341 N23341 0 diode
R23342 N23341 N23342 10
D23342 N23342 0 diode
R23343 N23342 N23343 10
D23343 N23343 0 diode
R23344 N23343 N23344 10
D23344 N23344 0 diode
R23345 N23344 N23345 10
D23345 N23345 0 diode
R23346 N23345 N23346 10
D23346 N23346 0 diode
R23347 N23346 N23347 10
D23347 N23347 0 diode
R23348 N23347 N23348 10
D23348 N23348 0 diode
R23349 N23348 N23349 10
D23349 N23349 0 diode
R23350 N23349 N23350 10
D23350 N23350 0 diode
R23351 N23350 N23351 10
D23351 N23351 0 diode
R23352 N23351 N23352 10
D23352 N23352 0 diode
R23353 N23352 N23353 10
D23353 N23353 0 diode
R23354 N23353 N23354 10
D23354 N23354 0 diode
R23355 N23354 N23355 10
D23355 N23355 0 diode
R23356 N23355 N23356 10
D23356 N23356 0 diode
R23357 N23356 N23357 10
D23357 N23357 0 diode
R23358 N23357 N23358 10
D23358 N23358 0 diode
R23359 N23358 N23359 10
D23359 N23359 0 diode
R23360 N23359 N23360 10
D23360 N23360 0 diode
R23361 N23360 N23361 10
D23361 N23361 0 diode
R23362 N23361 N23362 10
D23362 N23362 0 diode
R23363 N23362 N23363 10
D23363 N23363 0 diode
R23364 N23363 N23364 10
D23364 N23364 0 diode
R23365 N23364 N23365 10
D23365 N23365 0 diode
R23366 N23365 N23366 10
D23366 N23366 0 diode
R23367 N23366 N23367 10
D23367 N23367 0 diode
R23368 N23367 N23368 10
D23368 N23368 0 diode
R23369 N23368 N23369 10
D23369 N23369 0 diode
R23370 N23369 N23370 10
D23370 N23370 0 diode
R23371 N23370 N23371 10
D23371 N23371 0 diode
R23372 N23371 N23372 10
D23372 N23372 0 diode
R23373 N23372 N23373 10
D23373 N23373 0 diode
R23374 N23373 N23374 10
D23374 N23374 0 diode
R23375 N23374 N23375 10
D23375 N23375 0 diode
R23376 N23375 N23376 10
D23376 N23376 0 diode
R23377 N23376 N23377 10
D23377 N23377 0 diode
R23378 N23377 N23378 10
D23378 N23378 0 diode
R23379 N23378 N23379 10
D23379 N23379 0 diode
R23380 N23379 N23380 10
D23380 N23380 0 diode
R23381 N23380 N23381 10
D23381 N23381 0 diode
R23382 N23381 N23382 10
D23382 N23382 0 diode
R23383 N23382 N23383 10
D23383 N23383 0 diode
R23384 N23383 N23384 10
D23384 N23384 0 diode
R23385 N23384 N23385 10
D23385 N23385 0 diode
R23386 N23385 N23386 10
D23386 N23386 0 diode
R23387 N23386 N23387 10
D23387 N23387 0 diode
R23388 N23387 N23388 10
D23388 N23388 0 diode
R23389 N23388 N23389 10
D23389 N23389 0 diode
R23390 N23389 N23390 10
D23390 N23390 0 diode
R23391 N23390 N23391 10
D23391 N23391 0 diode
R23392 N23391 N23392 10
D23392 N23392 0 diode
R23393 N23392 N23393 10
D23393 N23393 0 diode
R23394 N23393 N23394 10
D23394 N23394 0 diode
R23395 N23394 N23395 10
D23395 N23395 0 diode
R23396 N23395 N23396 10
D23396 N23396 0 diode
R23397 N23396 N23397 10
D23397 N23397 0 diode
R23398 N23397 N23398 10
D23398 N23398 0 diode
R23399 N23398 N23399 10
D23399 N23399 0 diode
R23400 N23399 N23400 10
D23400 N23400 0 diode
R23401 N23400 N23401 10
D23401 N23401 0 diode
R23402 N23401 N23402 10
D23402 N23402 0 diode
R23403 N23402 N23403 10
D23403 N23403 0 diode
R23404 N23403 N23404 10
D23404 N23404 0 diode
R23405 N23404 N23405 10
D23405 N23405 0 diode
R23406 N23405 N23406 10
D23406 N23406 0 diode
R23407 N23406 N23407 10
D23407 N23407 0 diode
R23408 N23407 N23408 10
D23408 N23408 0 diode
R23409 N23408 N23409 10
D23409 N23409 0 diode
R23410 N23409 N23410 10
D23410 N23410 0 diode
R23411 N23410 N23411 10
D23411 N23411 0 diode
R23412 N23411 N23412 10
D23412 N23412 0 diode
R23413 N23412 N23413 10
D23413 N23413 0 diode
R23414 N23413 N23414 10
D23414 N23414 0 diode
R23415 N23414 N23415 10
D23415 N23415 0 diode
R23416 N23415 N23416 10
D23416 N23416 0 diode
R23417 N23416 N23417 10
D23417 N23417 0 diode
R23418 N23417 N23418 10
D23418 N23418 0 diode
R23419 N23418 N23419 10
D23419 N23419 0 diode
R23420 N23419 N23420 10
D23420 N23420 0 diode
R23421 N23420 N23421 10
D23421 N23421 0 diode
R23422 N23421 N23422 10
D23422 N23422 0 diode
R23423 N23422 N23423 10
D23423 N23423 0 diode
R23424 N23423 N23424 10
D23424 N23424 0 diode
R23425 N23424 N23425 10
D23425 N23425 0 diode
R23426 N23425 N23426 10
D23426 N23426 0 diode
R23427 N23426 N23427 10
D23427 N23427 0 diode
R23428 N23427 N23428 10
D23428 N23428 0 diode
R23429 N23428 N23429 10
D23429 N23429 0 diode
R23430 N23429 N23430 10
D23430 N23430 0 diode
R23431 N23430 N23431 10
D23431 N23431 0 diode
R23432 N23431 N23432 10
D23432 N23432 0 diode
R23433 N23432 N23433 10
D23433 N23433 0 diode
R23434 N23433 N23434 10
D23434 N23434 0 diode
R23435 N23434 N23435 10
D23435 N23435 0 diode
R23436 N23435 N23436 10
D23436 N23436 0 diode
R23437 N23436 N23437 10
D23437 N23437 0 diode
R23438 N23437 N23438 10
D23438 N23438 0 diode
R23439 N23438 N23439 10
D23439 N23439 0 diode
R23440 N23439 N23440 10
D23440 N23440 0 diode
R23441 N23440 N23441 10
D23441 N23441 0 diode
R23442 N23441 N23442 10
D23442 N23442 0 diode
R23443 N23442 N23443 10
D23443 N23443 0 diode
R23444 N23443 N23444 10
D23444 N23444 0 diode
R23445 N23444 N23445 10
D23445 N23445 0 diode
R23446 N23445 N23446 10
D23446 N23446 0 diode
R23447 N23446 N23447 10
D23447 N23447 0 diode
R23448 N23447 N23448 10
D23448 N23448 0 diode
R23449 N23448 N23449 10
D23449 N23449 0 diode
R23450 N23449 N23450 10
D23450 N23450 0 diode
R23451 N23450 N23451 10
D23451 N23451 0 diode
R23452 N23451 N23452 10
D23452 N23452 0 diode
R23453 N23452 N23453 10
D23453 N23453 0 diode
R23454 N23453 N23454 10
D23454 N23454 0 diode
R23455 N23454 N23455 10
D23455 N23455 0 diode
R23456 N23455 N23456 10
D23456 N23456 0 diode
R23457 N23456 N23457 10
D23457 N23457 0 diode
R23458 N23457 N23458 10
D23458 N23458 0 diode
R23459 N23458 N23459 10
D23459 N23459 0 diode
R23460 N23459 N23460 10
D23460 N23460 0 diode
R23461 N23460 N23461 10
D23461 N23461 0 diode
R23462 N23461 N23462 10
D23462 N23462 0 diode
R23463 N23462 N23463 10
D23463 N23463 0 diode
R23464 N23463 N23464 10
D23464 N23464 0 diode
R23465 N23464 N23465 10
D23465 N23465 0 diode
R23466 N23465 N23466 10
D23466 N23466 0 diode
R23467 N23466 N23467 10
D23467 N23467 0 diode
R23468 N23467 N23468 10
D23468 N23468 0 diode
R23469 N23468 N23469 10
D23469 N23469 0 diode
R23470 N23469 N23470 10
D23470 N23470 0 diode
R23471 N23470 N23471 10
D23471 N23471 0 diode
R23472 N23471 N23472 10
D23472 N23472 0 diode
R23473 N23472 N23473 10
D23473 N23473 0 diode
R23474 N23473 N23474 10
D23474 N23474 0 diode
R23475 N23474 N23475 10
D23475 N23475 0 diode
R23476 N23475 N23476 10
D23476 N23476 0 diode
R23477 N23476 N23477 10
D23477 N23477 0 diode
R23478 N23477 N23478 10
D23478 N23478 0 diode
R23479 N23478 N23479 10
D23479 N23479 0 diode
R23480 N23479 N23480 10
D23480 N23480 0 diode
R23481 N23480 N23481 10
D23481 N23481 0 diode
R23482 N23481 N23482 10
D23482 N23482 0 diode
R23483 N23482 N23483 10
D23483 N23483 0 diode
R23484 N23483 N23484 10
D23484 N23484 0 diode
R23485 N23484 N23485 10
D23485 N23485 0 diode
R23486 N23485 N23486 10
D23486 N23486 0 diode
R23487 N23486 N23487 10
D23487 N23487 0 diode
R23488 N23487 N23488 10
D23488 N23488 0 diode
R23489 N23488 N23489 10
D23489 N23489 0 diode
R23490 N23489 N23490 10
D23490 N23490 0 diode
R23491 N23490 N23491 10
D23491 N23491 0 diode
R23492 N23491 N23492 10
D23492 N23492 0 diode
R23493 N23492 N23493 10
D23493 N23493 0 diode
R23494 N23493 N23494 10
D23494 N23494 0 diode
R23495 N23494 N23495 10
D23495 N23495 0 diode
R23496 N23495 N23496 10
D23496 N23496 0 diode
R23497 N23496 N23497 10
D23497 N23497 0 diode
R23498 N23497 N23498 10
D23498 N23498 0 diode
R23499 N23498 N23499 10
D23499 N23499 0 diode
R23500 N23499 N23500 10
D23500 N23500 0 diode
R23501 N23500 N23501 10
D23501 N23501 0 diode
R23502 N23501 N23502 10
D23502 N23502 0 diode
R23503 N23502 N23503 10
D23503 N23503 0 diode
R23504 N23503 N23504 10
D23504 N23504 0 diode
R23505 N23504 N23505 10
D23505 N23505 0 diode
R23506 N23505 N23506 10
D23506 N23506 0 diode
R23507 N23506 N23507 10
D23507 N23507 0 diode
R23508 N23507 N23508 10
D23508 N23508 0 diode
R23509 N23508 N23509 10
D23509 N23509 0 diode
R23510 N23509 N23510 10
D23510 N23510 0 diode
R23511 N23510 N23511 10
D23511 N23511 0 diode
R23512 N23511 N23512 10
D23512 N23512 0 diode
R23513 N23512 N23513 10
D23513 N23513 0 diode
R23514 N23513 N23514 10
D23514 N23514 0 diode
R23515 N23514 N23515 10
D23515 N23515 0 diode
R23516 N23515 N23516 10
D23516 N23516 0 diode
R23517 N23516 N23517 10
D23517 N23517 0 diode
R23518 N23517 N23518 10
D23518 N23518 0 diode
R23519 N23518 N23519 10
D23519 N23519 0 diode
R23520 N23519 N23520 10
D23520 N23520 0 diode
R23521 N23520 N23521 10
D23521 N23521 0 diode
R23522 N23521 N23522 10
D23522 N23522 0 diode
R23523 N23522 N23523 10
D23523 N23523 0 diode
R23524 N23523 N23524 10
D23524 N23524 0 diode
R23525 N23524 N23525 10
D23525 N23525 0 diode
R23526 N23525 N23526 10
D23526 N23526 0 diode
R23527 N23526 N23527 10
D23527 N23527 0 diode
R23528 N23527 N23528 10
D23528 N23528 0 diode
R23529 N23528 N23529 10
D23529 N23529 0 diode
R23530 N23529 N23530 10
D23530 N23530 0 diode
R23531 N23530 N23531 10
D23531 N23531 0 diode
R23532 N23531 N23532 10
D23532 N23532 0 diode
R23533 N23532 N23533 10
D23533 N23533 0 diode
R23534 N23533 N23534 10
D23534 N23534 0 diode
R23535 N23534 N23535 10
D23535 N23535 0 diode
R23536 N23535 N23536 10
D23536 N23536 0 diode
R23537 N23536 N23537 10
D23537 N23537 0 diode
R23538 N23537 N23538 10
D23538 N23538 0 diode
R23539 N23538 N23539 10
D23539 N23539 0 diode
R23540 N23539 N23540 10
D23540 N23540 0 diode
R23541 N23540 N23541 10
D23541 N23541 0 diode
R23542 N23541 N23542 10
D23542 N23542 0 diode
R23543 N23542 N23543 10
D23543 N23543 0 diode
R23544 N23543 N23544 10
D23544 N23544 0 diode
R23545 N23544 N23545 10
D23545 N23545 0 diode
R23546 N23545 N23546 10
D23546 N23546 0 diode
R23547 N23546 N23547 10
D23547 N23547 0 diode
R23548 N23547 N23548 10
D23548 N23548 0 diode
R23549 N23548 N23549 10
D23549 N23549 0 diode
R23550 N23549 N23550 10
D23550 N23550 0 diode
R23551 N23550 N23551 10
D23551 N23551 0 diode
R23552 N23551 N23552 10
D23552 N23552 0 diode
R23553 N23552 N23553 10
D23553 N23553 0 diode
R23554 N23553 N23554 10
D23554 N23554 0 diode
R23555 N23554 N23555 10
D23555 N23555 0 diode
R23556 N23555 N23556 10
D23556 N23556 0 diode
R23557 N23556 N23557 10
D23557 N23557 0 diode
R23558 N23557 N23558 10
D23558 N23558 0 diode
R23559 N23558 N23559 10
D23559 N23559 0 diode
R23560 N23559 N23560 10
D23560 N23560 0 diode
R23561 N23560 N23561 10
D23561 N23561 0 diode
R23562 N23561 N23562 10
D23562 N23562 0 diode
R23563 N23562 N23563 10
D23563 N23563 0 diode
R23564 N23563 N23564 10
D23564 N23564 0 diode
R23565 N23564 N23565 10
D23565 N23565 0 diode
R23566 N23565 N23566 10
D23566 N23566 0 diode
R23567 N23566 N23567 10
D23567 N23567 0 diode
R23568 N23567 N23568 10
D23568 N23568 0 diode
R23569 N23568 N23569 10
D23569 N23569 0 diode
R23570 N23569 N23570 10
D23570 N23570 0 diode
R23571 N23570 N23571 10
D23571 N23571 0 diode
R23572 N23571 N23572 10
D23572 N23572 0 diode
R23573 N23572 N23573 10
D23573 N23573 0 diode
R23574 N23573 N23574 10
D23574 N23574 0 diode
R23575 N23574 N23575 10
D23575 N23575 0 diode
R23576 N23575 N23576 10
D23576 N23576 0 diode
R23577 N23576 N23577 10
D23577 N23577 0 diode
R23578 N23577 N23578 10
D23578 N23578 0 diode
R23579 N23578 N23579 10
D23579 N23579 0 diode
R23580 N23579 N23580 10
D23580 N23580 0 diode
R23581 N23580 N23581 10
D23581 N23581 0 diode
R23582 N23581 N23582 10
D23582 N23582 0 diode
R23583 N23582 N23583 10
D23583 N23583 0 diode
R23584 N23583 N23584 10
D23584 N23584 0 diode
R23585 N23584 N23585 10
D23585 N23585 0 diode
R23586 N23585 N23586 10
D23586 N23586 0 diode
R23587 N23586 N23587 10
D23587 N23587 0 diode
R23588 N23587 N23588 10
D23588 N23588 0 diode
R23589 N23588 N23589 10
D23589 N23589 0 diode
R23590 N23589 N23590 10
D23590 N23590 0 diode
R23591 N23590 N23591 10
D23591 N23591 0 diode
R23592 N23591 N23592 10
D23592 N23592 0 diode
R23593 N23592 N23593 10
D23593 N23593 0 diode
R23594 N23593 N23594 10
D23594 N23594 0 diode
R23595 N23594 N23595 10
D23595 N23595 0 diode
R23596 N23595 N23596 10
D23596 N23596 0 diode
R23597 N23596 N23597 10
D23597 N23597 0 diode
R23598 N23597 N23598 10
D23598 N23598 0 diode
R23599 N23598 N23599 10
D23599 N23599 0 diode
R23600 N23599 N23600 10
D23600 N23600 0 diode
R23601 N23600 N23601 10
D23601 N23601 0 diode
R23602 N23601 N23602 10
D23602 N23602 0 diode
R23603 N23602 N23603 10
D23603 N23603 0 diode
R23604 N23603 N23604 10
D23604 N23604 0 diode
R23605 N23604 N23605 10
D23605 N23605 0 diode
R23606 N23605 N23606 10
D23606 N23606 0 diode
R23607 N23606 N23607 10
D23607 N23607 0 diode
R23608 N23607 N23608 10
D23608 N23608 0 diode
R23609 N23608 N23609 10
D23609 N23609 0 diode
R23610 N23609 N23610 10
D23610 N23610 0 diode
R23611 N23610 N23611 10
D23611 N23611 0 diode
R23612 N23611 N23612 10
D23612 N23612 0 diode
R23613 N23612 N23613 10
D23613 N23613 0 diode
R23614 N23613 N23614 10
D23614 N23614 0 diode
R23615 N23614 N23615 10
D23615 N23615 0 diode
R23616 N23615 N23616 10
D23616 N23616 0 diode
R23617 N23616 N23617 10
D23617 N23617 0 diode
R23618 N23617 N23618 10
D23618 N23618 0 diode
R23619 N23618 N23619 10
D23619 N23619 0 diode
R23620 N23619 N23620 10
D23620 N23620 0 diode
R23621 N23620 N23621 10
D23621 N23621 0 diode
R23622 N23621 N23622 10
D23622 N23622 0 diode
R23623 N23622 N23623 10
D23623 N23623 0 diode
R23624 N23623 N23624 10
D23624 N23624 0 diode
R23625 N23624 N23625 10
D23625 N23625 0 diode
R23626 N23625 N23626 10
D23626 N23626 0 diode
R23627 N23626 N23627 10
D23627 N23627 0 diode
R23628 N23627 N23628 10
D23628 N23628 0 diode
R23629 N23628 N23629 10
D23629 N23629 0 diode
R23630 N23629 N23630 10
D23630 N23630 0 diode
R23631 N23630 N23631 10
D23631 N23631 0 diode
R23632 N23631 N23632 10
D23632 N23632 0 diode
R23633 N23632 N23633 10
D23633 N23633 0 diode
R23634 N23633 N23634 10
D23634 N23634 0 diode
R23635 N23634 N23635 10
D23635 N23635 0 diode
R23636 N23635 N23636 10
D23636 N23636 0 diode
R23637 N23636 N23637 10
D23637 N23637 0 diode
R23638 N23637 N23638 10
D23638 N23638 0 diode
R23639 N23638 N23639 10
D23639 N23639 0 diode
R23640 N23639 N23640 10
D23640 N23640 0 diode
R23641 N23640 N23641 10
D23641 N23641 0 diode
R23642 N23641 N23642 10
D23642 N23642 0 diode
R23643 N23642 N23643 10
D23643 N23643 0 diode
R23644 N23643 N23644 10
D23644 N23644 0 diode
R23645 N23644 N23645 10
D23645 N23645 0 diode
R23646 N23645 N23646 10
D23646 N23646 0 diode
R23647 N23646 N23647 10
D23647 N23647 0 diode
R23648 N23647 N23648 10
D23648 N23648 0 diode
R23649 N23648 N23649 10
D23649 N23649 0 diode
R23650 N23649 N23650 10
D23650 N23650 0 diode
R23651 N23650 N23651 10
D23651 N23651 0 diode
R23652 N23651 N23652 10
D23652 N23652 0 diode
R23653 N23652 N23653 10
D23653 N23653 0 diode
R23654 N23653 N23654 10
D23654 N23654 0 diode
R23655 N23654 N23655 10
D23655 N23655 0 diode
R23656 N23655 N23656 10
D23656 N23656 0 diode
R23657 N23656 N23657 10
D23657 N23657 0 diode
R23658 N23657 N23658 10
D23658 N23658 0 diode
R23659 N23658 N23659 10
D23659 N23659 0 diode
R23660 N23659 N23660 10
D23660 N23660 0 diode
R23661 N23660 N23661 10
D23661 N23661 0 diode
R23662 N23661 N23662 10
D23662 N23662 0 diode
R23663 N23662 N23663 10
D23663 N23663 0 diode
R23664 N23663 N23664 10
D23664 N23664 0 diode
R23665 N23664 N23665 10
D23665 N23665 0 diode
R23666 N23665 N23666 10
D23666 N23666 0 diode
R23667 N23666 N23667 10
D23667 N23667 0 diode
R23668 N23667 N23668 10
D23668 N23668 0 diode
R23669 N23668 N23669 10
D23669 N23669 0 diode
R23670 N23669 N23670 10
D23670 N23670 0 diode
R23671 N23670 N23671 10
D23671 N23671 0 diode
R23672 N23671 N23672 10
D23672 N23672 0 diode
R23673 N23672 N23673 10
D23673 N23673 0 diode
R23674 N23673 N23674 10
D23674 N23674 0 diode
R23675 N23674 N23675 10
D23675 N23675 0 diode
R23676 N23675 N23676 10
D23676 N23676 0 diode
R23677 N23676 N23677 10
D23677 N23677 0 diode
R23678 N23677 N23678 10
D23678 N23678 0 diode
R23679 N23678 N23679 10
D23679 N23679 0 diode
R23680 N23679 N23680 10
D23680 N23680 0 diode
R23681 N23680 N23681 10
D23681 N23681 0 diode
R23682 N23681 N23682 10
D23682 N23682 0 diode
R23683 N23682 N23683 10
D23683 N23683 0 diode
R23684 N23683 N23684 10
D23684 N23684 0 diode
R23685 N23684 N23685 10
D23685 N23685 0 diode
R23686 N23685 N23686 10
D23686 N23686 0 diode
R23687 N23686 N23687 10
D23687 N23687 0 diode
R23688 N23687 N23688 10
D23688 N23688 0 diode
R23689 N23688 N23689 10
D23689 N23689 0 diode
R23690 N23689 N23690 10
D23690 N23690 0 diode
R23691 N23690 N23691 10
D23691 N23691 0 diode
R23692 N23691 N23692 10
D23692 N23692 0 diode
R23693 N23692 N23693 10
D23693 N23693 0 diode
R23694 N23693 N23694 10
D23694 N23694 0 diode
R23695 N23694 N23695 10
D23695 N23695 0 diode
R23696 N23695 N23696 10
D23696 N23696 0 diode
R23697 N23696 N23697 10
D23697 N23697 0 diode
R23698 N23697 N23698 10
D23698 N23698 0 diode
R23699 N23698 N23699 10
D23699 N23699 0 diode
R23700 N23699 N23700 10
D23700 N23700 0 diode
R23701 N23700 N23701 10
D23701 N23701 0 diode
R23702 N23701 N23702 10
D23702 N23702 0 diode
R23703 N23702 N23703 10
D23703 N23703 0 diode
R23704 N23703 N23704 10
D23704 N23704 0 diode
R23705 N23704 N23705 10
D23705 N23705 0 diode
R23706 N23705 N23706 10
D23706 N23706 0 diode
R23707 N23706 N23707 10
D23707 N23707 0 diode
R23708 N23707 N23708 10
D23708 N23708 0 diode
R23709 N23708 N23709 10
D23709 N23709 0 diode
R23710 N23709 N23710 10
D23710 N23710 0 diode
R23711 N23710 N23711 10
D23711 N23711 0 diode
R23712 N23711 N23712 10
D23712 N23712 0 diode
R23713 N23712 N23713 10
D23713 N23713 0 diode
R23714 N23713 N23714 10
D23714 N23714 0 diode
R23715 N23714 N23715 10
D23715 N23715 0 diode
R23716 N23715 N23716 10
D23716 N23716 0 diode
R23717 N23716 N23717 10
D23717 N23717 0 diode
R23718 N23717 N23718 10
D23718 N23718 0 diode
R23719 N23718 N23719 10
D23719 N23719 0 diode
R23720 N23719 N23720 10
D23720 N23720 0 diode
R23721 N23720 N23721 10
D23721 N23721 0 diode
R23722 N23721 N23722 10
D23722 N23722 0 diode
R23723 N23722 N23723 10
D23723 N23723 0 diode
R23724 N23723 N23724 10
D23724 N23724 0 diode
R23725 N23724 N23725 10
D23725 N23725 0 diode
R23726 N23725 N23726 10
D23726 N23726 0 diode
R23727 N23726 N23727 10
D23727 N23727 0 diode
R23728 N23727 N23728 10
D23728 N23728 0 diode
R23729 N23728 N23729 10
D23729 N23729 0 diode
R23730 N23729 N23730 10
D23730 N23730 0 diode
R23731 N23730 N23731 10
D23731 N23731 0 diode
R23732 N23731 N23732 10
D23732 N23732 0 diode
R23733 N23732 N23733 10
D23733 N23733 0 diode
R23734 N23733 N23734 10
D23734 N23734 0 diode
R23735 N23734 N23735 10
D23735 N23735 0 diode
R23736 N23735 N23736 10
D23736 N23736 0 diode
R23737 N23736 N23737 10
D23737 N23737 0 diode
R23738 N23737 N23738 10
D23738 N23738 0 diode
R23739 N23738 N23739 10
D23739 N23739 0 diode
R23740 N23739 N23740 10
D23740 N23740 0 diode
R23741 N23740 N23741 10
D23741 N23741 0 diode
R23742 N23741 N23742 10
D23742 N23742 0 diode
R23743 N23742 N23743 10
D23743 N23743 0 diode
R23744 N23743 N23744 10
D23744 N23744 0 diode
R23745 N23744 N23745 10
D23745 N23745 0 diode
R23746 N23745 N23746 10
D23746 N23746 0 diode
R23747 N23746 N23747 10
D23747 N23747 0 diode
R23748 N23747 N23748 10
D23748 N23748 0 diode
R23749 N23748 N23749 10
D23749 N23749 0 diode
R23750 N23749 N23750 10
D23750 N23750 0 diode
R23751 N23750 N23751 10
D23751 N23751 0 diode
R23752 N23751 N23752 10
D23752 N23752 0 diode
R23753 N23752 N23753 10
D23753 N23753 0 diode
R23754 N23753 N23754 10
D23754 N23754 0 diode
R23755 N23754 N23755 10
D23755 N23755 0 diode
R23756 N23755 N23756 10
D23756 N23756 0 diode
R23757 N23756 N23757 10
D23757 N23757 0 diode
R23758 N23757 N23758 10
D23758 N23758 0 diode
R23759 N23758 N23759 10
D23759 N23759 0 diode
R23760 N23759 N23760 10
D23760 N23760 0 diode
R23761 N23760 N23761 10
D23761 N23761 0 diode
R23762 N23761 N23762 10
D23762 N23762 0 diode
R23763 N23762 N23763 10
D23763 N23763 0 diode
R23764 N23763 N23764 10
D23764 N23764 0 diode
R23765 N23764 N23765 10
D23765 N23765 0 diode
R23766 N23765 N23766 10
D23766 N23766 0 diode
R23767 N23766 N23767 10
D23767 N23767 0 diode
R23768 N23767 N23768 10
D23768 N23768 0 diode
R23769 N23768 N23769 10
D23769 N23769 0 diode
R23770 N23769 N23770 10
D23770 N23770 0 diode
R23771 N23770 N23771 10
D23771 N23771 0 diode
R23772 N23771 N23772 10
D23772 N23772 0 diode
R23773 N23772 N23773 10
D23773 N23773 0 diode
R23774 N23773 N23774 10
D23774 N23774 0 diode
R23775 N23774 N23775 10
D23775 N23775 0 diode
R23776 N23775 N23776 10
D23776 N23776 0 diode
R23777 N23776 N23777 10
D23777 N23777 0 diode
R23778 N23777 N23778 10
D23778 N23778 0 diode
R23779 N23778 N23779 10
D23779 N23779 0 diode
R23780 N23779 N23780 10
D23780 N23780 0 diode
R23781 N23780 N23781 10
D23781 N23781 0 diode
R23782 N23781 N23782 10
D23782 N23782 0 diode
R23783 N23782 N23783 10
D23783 N23783 0 diode
R23784 N23783 N23784 10
D23784 N23784 0 diode
R23785 N23784 N23785 10
D23785 N23785 0 diode
R23786 N23785 N23786 10
D23786 N23786 0 diode
R23787 N23786 N23787 10
D23787 N23787 0 diode
R23788 N23787 N23788 10
D23788 N23788 0 diode
R23789 N23788 N23789 10
D23789 N23789 0 diode
R23790 N23789 N23790 10
D23790 N23790 0 diode
R23791 N23790 N23791 10
D23791 N23791 0 diode
R23792 N23791 N23792 10
D23792 N23792 0 diode
R23793 N23792 N23793 10
D23793 N23793 0 diode
R23794 N23793 N23794 10
D23794 N23794 0 diode
R23795 N23794 N23795 10
D23795 N23795 0 diode
R23796 N23795 N23796 10
D23796 N23796 0 diode
R23797 N23796 N23797 10
D23797 N23797 0 diode
R23798 N23797 N23798 10
D23798 N23798 0 diode
R23799 N23798 N23799 10
D23799 N23799 0 diode
R23800 N23799 N23800 10
D23800 N23800 0 diode
R23801 N23800 N23801 10
D23801 N23801 0 diode
R23802 N23801 N23802 10
D23802 N23802 0 diode
R23803 N23802 N23803 10
D23803 N23803 0 diode
R23804 N23803 N23804 10
D23804 N23804 0 diode
R23805 N23804 N23805 10
D23805 N23805 0 diode
R23806 N23805 N23806 10
D23806 N23806 0 diode
R23807 N23806 N23807 10
D23807 N23807 0 diode
R23808 N23807 N23808 10
D23808 N23808 0 diode
R23809 N23808 N23809 10
D23809 N23809 0 diode
R23810 N23809 N23810 10
D23810 N23810 0 diode
R23811 N23810 N23811 10
D23811 N23811 0 diode
R23812 N23811 N23812 10
D23812 N23812 0 diode
R23813 N23812 N23813 10
D23813 N23813 0 diode
R23814 N23813 N23814 10
D23814 N23814 0 diode
R23815 N23814 N23815 10
D23815 N23815 0 diode
R23816 N23815 N23816 10
D23816 N23816 0 diode
R23817 N23816 N23817 10
D23817 N23817 0 diode
R23818 N23817 N23818 10
D23818 N23818 0 diode
R23819 N23818 N23819 10
D23819 N23819 0 diode
R23820 N23819 N23820 10
D23820 N23820 0 diode
R23821 N23820 N23821 10
D23821 N23821 0 diode
R23822 N23821 N23822 10
D23822 N23822 0 diode
R23823 N23822 N23823 10
D23823 N23823 0 diode
R23824 N23823 N23824 10
D23824 N23824 0 diode
R23825 N23824 N23825 10
D23825 N23825 0 diode
R23826 N23825 N23826 10
D23826 N23826 0 diode
R23827 N23826 N23827 10
D23827 N23827 0 diode
R23828 N23827 N23828 10
D23828 N23828 0 diode
R23829 N23828 N23829 10
D23829 N23829 0 diode
R23830 N23829 N23830 10
D23830 N23830 0 diode
R23831 N23830 N23831 10
D23831 N23831 0 diode
R23832 N23831 N23832 10
D23832 N23832 0 diode
R23833 N23832 N23833 10
D23833 N23833 0 diode
R23834 N23833 N23834 10
D23834 N23834 0 diode
R23835 N23834 N23835 10
D23835 N23835 0 diode
R23836 N23835 N23836 10
D23836 N23836 0 diode
R23837 N23836 N23837 10
D23837 N23837 0 diode
R23838 N23837 N23838 10
D23838 N23838 0 diode
R23839 N23838 N23839 10
D23839 N23839 0 diode
R23840 N23839 N23840 10
D23840 N23840 0 diode
R23841 N23840 N23841 10
D23841 N23841 0 diode
R23842 N23841 N23842 10
D23842 N23842 0 diode
R23843 N23842 N23843 10
D23843 N23843 0 diode
R23844 N23843 N23844 10
D23844 N23844 0 diode
R23845 N23844 N23845 10
D23845 N23845 0 diode
R23846 N23845 N23846 10
D23846 N23846 0 diode
R23847 N23846 N23847 10
D23847 N23847 0 diode
R23848 N23847 N23848 10
D23848 N23848 0 diode
R23849 N23848 N23849 10
D23849 N23849 0 diode
R23850 N23849 N23850 10
D23850 N23850 0 diode
R23851 N23850 N23851 10
D23851 N23851 0 diode
R23852 N23851 N23852 10
D23852 N23852 0 diode
R23853 N23852 N23853 10
D23853 N23853 0 diode
R23854 N23853 N23854 10
D23854 N23854 0 diode
R23855 N23854 N23855 10
D23855 N23855 0 diode
R23856 N23855 N23856 10
D23856 N23856 0 diode
R23857 N23856 N23857 10
D23857 N23857 0 diode
R23858 N23857 N23858 10
D23858 N23858 0 diode
R23859 N23858 N23859 10
D23859 N23859 0 diode
R23860 N23859 N23860 10
D23860 N23860 0 diode
R23861 N23860 N23861 10
D23861 N23861 0 diode
R23862 N23861 N23862 10
D23862 N23862 0 diode
R23863 N23862 N23863 10
D23863 N23863 0 diode
R23864 N23863 N23864 10
D23864 N23864 0 diode
R23865 N23864 N23865 10
D23865 N23865 0 diode
R23866 N23865 N23866 10
D23866 N23866 0 diode
R23867 N23866 N23867 10
D23867 N23867 0 diode
R23868 N23867 N23868 10
D23868 N23868 0 diode
R23869 N23868 N23869 10
D23869 N23869 0 diode
R23870 N23869 N23870 10
D23870 N23870 0 diode
R23871 N23870 N23871 10
D23871 N23871 0 diode
R23872 N23871 N23872 10
D23872 N23872 0 diode
R23873 N23872 N23873 10
D23873 N23873 0 diode
R23874 N23873 N23874 10
D23874 N23874 0 diode
R23875 N23874 N23875 10
D23875 N23875 0 diode
R23876 N23875 N23876 10
D23876 N23876 0 diode
R23877 N23876 N23877 10
D23877 N23877 0 diode
R23878 N23877 N23878 10
D23878 N23878 0 diode
R23879 N23878 N23879 10
D23879 N23879 0 diode
R23880 N23879 N23880 10
D23880 N23880 0 diode
R23881 N23880 N23881 10
D23881 N23881 0 diode
R23882 N23881 N23882 10
D23882 N23882 0 diode
R23883 N23882 N23883 10
D23883 N23883 0 diode
R23884 N23883 N23884 10
D23884 N23884 0 diode
R23885 N23884 N23885 10
D23885 N23885 0 diode
R23886 N23885 N23886 10
D23886 N23886 0 diode
R23887 N23886 N23887 10
D23887 N23887 0 diode
R23888 N23887 N23888 10
D23888 N23888 0 diode
R23889 N23888 N23889 10
D23889 N23889 0 diode
R23890 N23889 N23890 10
D23890 N23890 0 diode
R23891 N23890 N23891 10
D23891 N23891 0 diode
R23892 N23891 N23892 10
D23892 N23892 0 diode
R23893 N23892 N23893 10
D23893 N23893 0 diode
R23894 N23893 N23894 10
D23894 N23894 0 diode
R23895 N23894 N23895 10
D23895 N23895 0 diode
R23896 N23895 N23896 10
D23896 N23896 0 diode
R23897 N23896 N23897 10
D23897 N23897 0 diode
R23898 N23897 N23898 10
D23898 N23898 0 diode
R23899 N23898 N23899 10
D23899 N23899 0 diode
R23900 N23899 N23900 10
D23900 N23900 0 diode
R23901 N23900 N23901 10
D23901 N23901 0 diode
R23902 N23901 N23902 10
D23902 N23902 0 diode
R23903 N23902 N23903 10
D23903 N23903 0 diode
R23904 N23903 N23904 10
D23904 N23904 0 diode
R23905 N23904 N23905 10
D23905 N23905 0 diode
R23906 N23905 N23906 10
D23906 N23906 0 diode
R23907 N23906 N23907 10
D23907 N23907 0 diode
R23908 N23907 N23908 10
D23908 N23908 0 diode
R23909 N23908 N23909 10
D23909 N23909 0 diode
R23910 N23909 N23910 10
D23910 N23910 0 diode
R23911 N23910 N23911 10
D23911 N23911 0 diode
R23912 N23911 N23912 10
D23912 N23912 0 diode
R23913 N23912 N23913 10
D23913 N23913 0 diode
R23914 N23913 N23914 10
D23914 N23914 0 diode
R23915 N23914 N23915 10
D23915 N23915 0 diode
R23916 N23915 N23916 10
D23916 N23916 0 diode
R23917 N23916 N23917 10
D23917 N23917 0 diode
R23918 N23917 N23918 10
D23918 N23918 0 diode
R23919 N23918 N23919 10
D23919 N23919 0 diode
R23920 N23919 N23920 10
D23920 N23920 0 diode
R23921 N23920 N23921 10
D23921 N23921 0 diode
R23922 N23921 N23922 10
D23922 N23922 0 diode
R23923 N23922 N23923 10
D23923 N23923 0 diode
R23924 N23923 N23924 10
D23924 N23924 0 diode
R23925 N23924 N23925 10
D23925 N23925 0 diode
R23926 N23925 N23926 10
D23926 N23926 0 diode
R23927 N23926 N23927 10
D23927 N23927 0 diode
R23928 N23927 N23928 10
D23928 N23928 0 diode
R23929 N23928 N23929 10
D23929 N23929 0 diode
R23930 N23929 N23930 10
D23930 N23930 0 diode
R23931 N23930 N23931 10
D23931 N23931 0 diode
R23932 N23931 N23932 10
D23932 N23932 0 diode
R23933 N23932 N23933 10
D23933 N23933 0 diode
R23934 N23933 N23934 10
D23934 N23934 0 diode
R23935 N23934 N23935 10
D23935 N23935 0 diode
R23936 N23935 N23936 10
D23936 N23936 0 diode
R23937 N23936 N23937 10
D23937 N23937 0 diode
R23938 N23937 N23938 10
D23938 N23938 0 diode
R23939 N23938 N23939 10
D23939 N23939 0 diode
R23940 N23939 N23940 10
D23940 N23940 0 diode
R23941 N23940 N23941 10
D23941 N23941 0 diode
R23942 N23941 N23942 10
D23942 N23942 0 diode
R23943 N23942 N23943 10
D23943 N23943 0 diode
R23944 N23943 N23944 10
D23944 N23944 0 diode
R23945 N23944 N23945 10
D23945 N23945 0 diode
R23946 N23945 N23946 10
D23946 N23946 0 diode
R23947 N23946 N23947 10
D23947 N23947 0 diode
R23948 N23947 N23948 10
D23948 N23948 0 diode
R23949 N23948 N23949 10
D23949 N23949 0 diode
R23950 N23949 N23950 10
D23950 N23950 0 diode
R23951 N23950 N23951 10
D23951 N23951 0 diode
R23952 N23951 N23952 10
D23952 N23952 0 diode
R23953 N23952 N23953 10
D23953 N23953 0 diode
R23954 N23953 N23954 10
D23954 N23954 0 diode
R23955 N23954 N23955 10
D23955 N23955 0 diode
R23956 N23955 N23956 10
D23956 N23956 0 diode
R23957 N23956 N23957 10
D23957 N23957 0 diode
R23958 N23957 N23958 10
D23958 N23958 0 diode
R23959 N23958 N23959 10
D23959 N23959 0 diode
R23960 N23959 N23960 10
D23960 N23960 0 diode
R23961 N23960 N23961 10
D23961 N23961 0 diode
R23962 N23961 N23962 10
D23962 N23962 0 diode
R23963 N23962 N23963 10
D23963 N23963 0 diode
R23964 N23963 N23964 10
D23964 N23964 0 diode
R23965 N23964 N23965 10
D23965 N23965 0 diode
R23966 N23965 N23966 10
D23966 N23966 0 diode
R23967 N23966 N23967 10
D23967 N23967 0 diode
R23968 N23967 N23968 10
D23968 N23968 0 diode
R23969 N23968 N23969 10
D23969 N23969 0 diode
R23970 N23969 N23970 10
D23970 N23970 0 diode
R23971 N23970 N23971 10
D23971 N23971 0 diode
R23972 N23971 N23972 10
D23972 N23972 0 diode
R23973 N23972 N23973 10
D23973 N23973 0 diode
R23974 N23973 N23974 10
D23974 N23974 0 diode
R23975 N23974 N23975 10
D23975 N23975 0 diode
R23976 N23975 N23976 10
D23976 N23976 0 diode
R23977 N23976 N23977 10
D23977 N23977 0 diode
R23978 N23977 N23978 10
D23978 N23978 0 diode
R23979 N23978 N23979 10
D23979 N23979 0 diode
R23980 N23979 N23980 10
D23980 N23980 0 diode
R23981 N23980 N23981 10
D23981 N23981 0 diode
R23982 N23981 N23982 10
D23982 N23982 0 diode
R23983 N23982 N23983 10
D23983 N23983 0 diode
R23984 N23983 N23984 10
D23984 N23984 0 diode
R23985 N23984 N23985 10
D23985 N23985 0 diode
R23986 N23985 N23986 10
D23986 N23986 0 diode
R23987 N23986 N23987 10
D23987 N23987 0 diode
R23988 N23987 N23988 10
D23988 N23988 0 diode
R23989 N23988 N23989 10
D23989 N23989 0 diode
R23990 N23989 N23990 10
D23990 N23990 0 diode
R23991 N23990 N23991 10
D23991 N23991 0 diode
R23992 N23991 N23992 10
D23992 N23992 0 diode
R23993 N23992 N23993 10
D23993 N23993 0 diode
R23994 N23993 N23994 10
D23994 N23994 0 diode
R23995 N23994 N23995 10
D23995 N23995 0 diode
R23996 N23995 N23996 10
D23996 N23996 0 diode
R23997 N23996 N23997 10
D23997 N23997 0 diode
R23998 N23997 N23998 10
D23998 N23998 0 diode
R23999 N23998 N23999 10
D23999 N23999 0 diode
R24000 N23999 N24000 10
D24000 N24000 0 diode
R24001 N24000 N24001 10
D24001 N24001 0 diode
R24002 N24001 N24002 10
D24002 N24002 0 diode
R24003 N24002 N24003 10
D24003 N24003 0 diode
R24004 N24003 N24004 10
D24004 N24004 0 diode
R24005 N24004 N24005 10
D24005 N24005 0 diode
R24006 N24005 N24006 10
D24006 N24006 0 diode
R24007 N24006 N24007 10
D24007 N24007 0 diode
R24008 N24007 N24008 10
D24008 N24008 0 diode
R24009 N24008 N24009 10
D24009 N24009 0 diode
R24010 N24009 N24010 10
D24010 N24010 0 diode
R24011 N24010 N24011 10
D24011 N24011 0 diode
R24012 N24011 N24012 10
D24012 N24012 0 diode
R24013 N24012 N24013 10
D24013 N24013 0 diode
R24014 N24013 N24014 10
D24014 N24014 0 diode
R24015 N24014 N24015 10
D24015 N24015 0 diode
R24016 N24015 N24016 10
D24016 N24016 0 diode
R24017 N24016 N24017 10
D24017 N24017 0 diode
R24018 N24017 N24018 10
D24018 N24018 0 diode
R24019 N24018 N24019 10
D24019 N24019 0 diode
R24020 N24019 N24020 10
D24020 N24020 0 diode
R24021 N24020 N24021 10
D24021 N24021 0 diode
R24022 N24021 N24022 10
D24022 N24022 0 diode
R24023 N24022 N24023 10
D24023 N24023 0 diode
R24024 N24023 N24024 10
D24024 N24024 0 diode
R24025 N24024 N24025 10
D24025 N24025 0 diode
R24026 N24025 N24026 10
D24026 N24026 0 diode
R24027 N24026 N24027 10
D24027 N24027 0 diode
R24028 N24027 N24028 10
D24028 N24028 0 diode
R24029 N24028 N24029 10
D24029 N24029 0 diode
R24030 N24029 N24030 10
D24030 N24030 0 diode
R24031 N24030 N24031 10
D24031 N24031 0 diode
R24032 N24031 N24032 10
D24032 N24032 0 diode
R24033 N24032 N24033 10
D24033 N24033 0 diode
R24034 N24033 N24034 10
D24034 N24034 0 diode
R24035 N24034 N24035 10
D24035 N24035 0 diode
R24036 N24035 N24036 10
D24036 N24036 0 diode
R24037 N24036 N24037 10
D24037 N24037 0 diode
R24038 N24037 N24038 10
D24038 N24038 0 diode
R24039 N24038 N24039 10
D24039 N24039 0 diode
R24040 N24039 N24040 10
D24040 N24040 0 diode
R24041 N24040 N24041 10
D24041 N24041 0 diode
R24042 N24041 N24042 10
D24042 N24042 0 diode
R24043 N24042 N24043 10
D24043 N24043 0 diode
R24044 N24043 N24044 10
D24044 N24044 0 diode
R24045 N24044 N24045 10
D24045 N24045 0 diode
R24046 N24045 N24046 10
D24046 N24046 0 diode
R24047 N24046 N24047 10
D24047 N24047 0 diode
R24048 N24047 N24048 10
D24048 N24048 0 diode
R24049 N24048 N24049 10
D24049 N24049 0 diode
R24050 N24049 N24050 10
D24050 N24050 0 diode
R24051 N24050 N24051 10
D24051 N24051 0 diode
R24052 N24051 N24052 10
D24052 N24052 0 diode
R24053 N24052 N24053 10
D24053 N24053 0 diode
R24054 N24053 N24054 10
D24054 N24054 0 diode
R24055 N24054 N24055 10
D24055 N24055 0 diode
R24056 N24055 N24056 10
D24056 N24056 0 diode
R24057 N24056 N24057 10
D24057 N24057 0 diode
R24058 N24057 N24058 10
D24058 N24058 0 diode
R24059 N24058 N24059 10
D24059 N24059 0 diode
R24060 N24059 N24060 10
D24060 N24060 0 diode
R24061 N24060 N24061 10
D24061 N24061 0 diode
R24062 N24061 N24062 10
D24062 N24062 0 diode
R24063 N24062 N24063 10
D24063 N24063 0 diode
R24064 N24063 N24064 10
D24064 N24064 0 diode
R24065 N24064 N24065 10
D24065 N24065 0 diode
R24066 N24065 N24066 10
D24066 N24066 0 diode
R24067 N24066 N24067 10
D24067 N24067 0 diode
R24068 N24067 N24068 10
D24068 N24068 0 diode
R24069 N24068 N24069 10
D24069 N24069 0 diode
R24070 N24069 N24070 10
D24070 N24070 0 diode
R24071 N24070 N24071 10
D24071 N24071 0 diode
R24072 N24071 N24072 10
D24072 N24072 0 diode
R24073 N24072 N24073 10
D24073 N24073 0 diode
R24074 N24073 N24074 10
D24074 N24074 0 diode
R24075 N24074 N24075 10
D24075 N24075 0 diode
R24076 N24075 N24076 10
D24076 N24076 0 diode
R24077 N24076 N24077 10
D24077 N24077 0 diode
R24078 N24077 N24078 10
D24078 N24078 0 diode
R24079 N24078 N24079 10
D24079 N24079 0 diode
R24080 N24079 N24080 10
D24080 N24080 0 diode
R24081 N24080 N24081 10
D24081 N24081 0 diode
R24082 N24081 N24082 10
D24082 N24082 0 diode
R24083 N24082 N24083 10
D24083 N24083 0 diode
R24084 N24083 N24084 10
D24084 N24084 0 diode
R24085 N24084 N24085 10
D24085 N24085 0 diode
R24086 N24085 N24086 10
D24086 N24086 0 diode
R24087 N24086 N24087 10
D24087 N24087 0 diode
R24088 N24087 N24088 10
D24088 N24088 0 diode
R24089 N24088 N24089 10
D24089 N24089 0 diode
R24090 N24089 N24090 10
D24090 N24090 0 diode
R24091 N24090 N24091 10
D24091 N24091 0 diode
R24092 N24091 N24092 10
D24092 N24092 0 diode
R24093 N24092 N24093 10
D24093 N24093 0 diode
R24094 N24093 N24094 10
D24094 N24094 0 diode
R24095 N24094 N24095 10
D24095 N24095 0 diode
R24096 N24095 N24096 10
D24096 N24096 0 diode
R24097 N24096 N24097 10
D24097 N24097 0 diode
R24098 N24097 N24098 10
D24098 N24098 0 diode
R24099 N24098 N24099 10
D24099 N24099 0 diode
R24100 N24099 N24100 10
D24100 N24100 0 diode
R24101 N24100 N24101 10
D24101 N24101 0 diode
R24102 N24101 N24102 10
D24102 N24102 0 diode
R24103 N24102 N24103 10
D24103 N24103 0 diode
R24104 N24103 N24104 10
D24104 N24104 0 diode
R24105 N24104 N24105 10
D24105 N24105 0 diode
R24106 N24105 N24106 10
D24106 N24106 0 diode
R24107 N24106 N24107 10
D24107 N24107 0 diode
R24108 N24107 N24108 10
D24108 N24108 0 diode
R24109 N24108 N24109 10
D24109 N24109 0 diode
R24110 N24109 N24110 10
D24110 N24110 0 diode
R24111 N24110 N24111 10
D24111 N24111 0 diode
R24112 N24111 N24112 10
D24112 N24112 0 diode
R24113 N24112 N24113 10
D24113 N24113 0 diode
R24114 N24113 N24114 10
D24114 N24114 0 diode
R24115 N24114 N24115 10
D24115 N24115 0 diode
R24116 N24115 N24116 10
D24116 N24116 0 diode
R24117 N24116 N24117 10
D24117 N24117 0 diode
R24118 N24117 N24118 10
D24118 N24118 0 diode
R24119 N24118 N24119 10
D24119 N24119 0 diode
R24120 N24119 N24120 10
D24120 N24120 0 diode
R24121 N24120 N24121 10
D24121 N24121 0 diode
R24122 N24121 N24122 10
D24122 N24122 0 diode
R24123 N24122 N24123 10
D24123 N24123 0 diode
R24124 N24123 N24124 10
D24124 N24124 0 diode
R24125 N24124 N24125 10
D24125 N24125 0 diode
R24126 N24125 N24126 10
D24126 N24126 0 diode
R24127 N24126 N24127 10
D24127 N24127 0 diode
R24128 N24127 N24128 10
D24128 N24128 0 diode
R24129 N24128 N24129 10
D24129 N24129 0 diode
R24130 N24129 N24130 10
D24130 N24130 0 diode
R24131 N24130 N24131 10
D24131 N24131 0 diode
R24132 N24131 N24132 10
D24132 N24132 0 diode
R24133 N24132 N24133 10
D24133 N24133 0 diode
R24134 N24133 N24134 10
D24134 N24134 0 diode
R24135 N24134 N24135 10
D24135 N24135 0 diode
R24136 N24135 N24136 10
D24136 N24136 0 diode
R24137 N24136 N24137 10
D24137 N24137 0 diode
R24138 N24137 N24138 10
D24138 N24138 0 diode
R24139 N24138 N24139 10
D24139 N24139 0 diode
R24140 N24139 N24140 10
D24140 N24140 0 diode
R24141 N24140 N24141 10
D24141 N24141 0 diode
R24142 N24141 N24142 10
D24142 N24142 0 diode
R24143 N24142 N24143 10
D24143 N24143 0 diode
R24144 N24143 N24144 10
D24144 N24144 0 diode
R24145 N24144 N24145 10
D24145 N24145 0 diode
R24146 N24145 N24146 10
D24146 N24146 0 diode
R24147 N24146 N24147 10
D24147 N24147 0 diode
R24148 N24147 N24148 10
D24148 N24148 0 diode
R24149 N24148 N24149 10
D24149 N24149 0 diode
R24150 N24149 N24150 10
D24150 N24150 0 diode
R24151 N24150 N24151 10
D24151 N24151 0 diode
R24152 N24151 N24152 10
D24152 N24152 0 diode
R24153 N24152 N24153 10
D24153 N24153 0 diode
R24154 N24153 N24154 10
D24154 N24154 0 diode
R24155 N24154 N24155 10
D24155 N24155 0 diode
R24156 N24155 N24156 10
D24156 N24156 0 diode
R24157 N24156 N24157 10
D24157 N24157 0 diode
R24158 N24157 N24158 10
D24158 N24158 0 diode
R24159 N24158 N24159 10
D24159 N24159 0 diode
R24160 N24159 N24160 10
D24160 N24160 0 diode
R24161 N24160 N24161 10
D24161 N24161 0 diode
R24162 N24161 N24162 10
D24162 N24162 0 diode
R24163 N24162 N24163 10
D24163 N24163 0 diode
R24164 N24163 N24164 10
D24164 N24164 0 diode
R24165 N24164 N24165 10
D24165 N24165 0 diode
R24166 N24165 N24166 10
D24166 N24166 0 diode
R24167 N24166 N24167 10
D24167 N24167 0 diode
R24168 N24167 N24168 10
D24168 N24168 0 diode
R24169 N24168 N24169 10
D24169 N24169 0 diode
R24170 N24169 N24170 10
D24170 N24170 0 diode
R24171 N24170 N24171 10
D24171 N24171 0 diode
R24172 N24171 N24172 10
D24172 N24172 0 diode
R24173 N24172 N24173 10
D24173 N24173 0 diode
R24174 N24173 N24174 10
D24174 N24174 0 diode
R24175 N24174 N24175 10
D24175 N24175 0 diode
R24176 N24175 N24176 10
D24176 N24176 0 diode
R24177 N24176 N24177 10
D24177 N24177 0 diode
R24178 N24177 N24178 10
D24178 N24178 0 diode
R24179 N24178 N24179 10
D24179 N24179 0 diode
R24180 N24179 N24180 10
D24180 N24180 0 diode
R24181 N24180 N24181 10
D24181 N24181 0 diode
R24182 N24181 N24182 10
D24182 N24182 0 diode
R24183 N24182 N24183 10
D24183 N24183 0 diode
R24184 N24183 N24184 10
D24184 N24184 0 diode
R24185 N24184 N24185 10
D24185 N24185 0 diode
R24186 N24185 N24186 10
D24186 N24186 0 diode
R24187 N24186 N24187 10
D24187 N24187 0 diode
R24188 N24187 N24188 10
D24188 N24188 0 diode
R24189 N24188 N24189 10
D24189 N24189 0 diode
R24190 N24189 N24190 10
D24190 N24190 0 diode
R24191 N24190 N24191 10
D24191 N24191 0 diode
R24192 N24191 N24192 10
D24192 N24192 0 diode
R24193 N24192 N24193 10
D24193 N24193 0 diode
R24194 N24193 N24194 10
D24194 N24194 0 diode
R24195 N24194 N24195 10
D24195 N24195 0 diode
R24196 N24195 N24196 10
D24196 N24196 0 diode
R24197 N24196 N24197 10
D24197 N24197 0 diode
R24198 N24197 N24198 10
D24198 N24198 0 diode
R24199 N24198 N24199 10
D24199 N24199 0 diode
R24200 N24199 N24200 10
D24200 N24200 0 diode
R24201 N24200 N24201 10
D24201 N24201 0 diode
R24202 N24201 N24202 10
D24202 N24202 0 diode
R24203 N24202 N24203 10
D24203 N24203 0 diode
R24204 N24203 N24204 10
D24204 N24204 0 diode
R24205 N24204 N24205 10
D24205 N24205 0 diode
R24206 N24205 N24206 10
D24206 N24206 0 diode
R24207 N24206 N24207 10
D24207 N24207 0 diode
R24208 N24207 N24208 10
D24208 N24208 0 diode
R24209 N24208 N24209 10
D24209 N24209 0 diode
R24210 N24209 N24210 10
D24210 N24210 0 diode
R24211 N24210 N24211 10
D24211 N24211 0 diode
R24212 N24211 N24212 10
D24212 N24212 0 diode
R24213 N24212 N24213 10
D24213 N24213 0 diode
R24214 N24213 N24214 10
D24214 N24214 0 diode
R24215 N24214 N24215 10
D24215 N24215 0 diode
R24216 N24215 N24216 10
D24216 N24216 0 diode
R24217 N24216 N24217 10
D24217 N24217 0 diode
R24218 N24217 N24218 10
D24218 N24218 0 diode
R24219 N24218 N24219 10
D24219 N24219 0 diode
R24220 N24219 N24220 10
D24220 N24220 0 diode
R24221 N24220 N24221 10
D24221 N24221 0 diode
R24222 N24221 N24222 10
D24222 N24222 0 diode
R24223 N24222 N24223 10
D24223 N24223 0 diode
R24224 N24223 N24224 10
D24224 N24224 0 diode
R24225 N24224 N24225 10
D24225 N24225 0 diode
R24226 N24225 N24226 10
D24226 N24226 0 diode
R24227 N24226 N24227 10
D24227 N24227 0 diode
R24228 N24227 N24228 10
D24228 N24228 0 diode
R24229 N24228 N24229 10
D24229 N24229 0 diode
R24230 N24229 N24230 10
D24230 N24230 0 diode
R24231 N24230 N24231 10
D24231 N24231 0 diode
R24232 N24231 N24232 10
D24232 N24232 0 diode
R24233 N24232 N24233 10
D24233 N24233 0 diode
R24234 N24233 N24234 10
D24234 N24234 0 diode
R24235 N24234 N24235 10
D24235 N24235 0 diode
R24236 N24235 N24236 10
D24236 N24236 0 diode
R24237 N24236 N24237 10
D24237 N24237 0 diode
R24238 N24237 N24238 10
D24238 N24238 0 diode
R24239 N24238 N24239 10
D24239 N24239 0 diode
R24240 N24239 N24240 10
D24240 N24240 0 diode
R24241 N24240 N24241 10
D24241 N24241 0 diode
R24242 N24241 N24242 10
D24242 N24242 0 diode
R24243 N24242 N24243 10
D24243 N24243 0 diode
R24244 N24243 N24244 10
D24244 N24244 0 diode
R24245 N24244 N24245 10
D24245 N24245 0 diode
R24246 N24245 N24246 10
D24246 N24246 0 diode
R24247 N24246 N24247 10
D24247 N24247 0 diode
R24248 N24247 N24248 10
D24248 N24248 0 diode
R24249 N24248 N24249 10
D24249 N24249 0 diode
R24250 N24249 N24250 10
D24250 N24250 0 diode
R24251 N24250 N24251 10
D24251 N24251 0 diode
R24252 N24251 N24252 10
D24252 N24252 0 diode
R24253 N24252 N24253 10
D24253 N24253 0 diode
R24254 N24253 N24254 10
D24254 N24254 0 diode
R24255 N24254 N24255 10
D24255 N24255 0 diode
R24256 N24255 N24256 10
D24256 N24256 0 diode
R24257 N24256 N24257 10
D24257 N24257 0 diode
R24258 N24257 N24258 10
D24258 N24258 0 diode
R24259 N24258 N24259 10
D24259 N24259 0 diode
R24260 N24259 N24260 10
D24260 N24260 0 diode
R24261 N24260 N24261 10
D24261 N24261 0 diode
R24262 N24261 N24262 10
D24262 N24262 0 diode
R24263 N24262 N24263 10
D24263 N24263 0 diode
R24264 N24263 N24264 10
D24264 N24264 0 diode
R24265 N24264 N24265 10
D24265 N24265 0 diode
R24266 N24265 N24266 10
D24266 N24266 0 diode
R24267 N24266 N24267 10
D24267 N24267 0 diode
R24268 N24267 N24268 10
D24268 N24268 0 diode
R24269 N24268 N24269 10
D24269 N24269 0 diode
R24270 N24269 N24270 10
D24270 N24270 0 diode
R24271 N24270 N24271 10
D24271 N24271 0 diode
R24272 N24271 N24272 10
D24272 N24272 0 diode
R24273 N24272 N24273 10
D24273 N24273 0 diode
R24274 N24273 N24274 10
D24274 N24274 0 diode
R24275 N24274 N24275 10
D24275 N24275 0 diode
R24276 N24275 N24276 10
D24276 N24276 0 diode
R24277 N24276 N24277 10
D24277 N24277 0 diode
R24278 N24277 N24278 10
D24278 N24278 0 diode
R24279 N24278 N24279 10
D24279 N24279 0 diode
R24280 N24279 N24280 10
D24280 N24280 0 diode
R24281 N24280 N24281 10
D24281 N24281 0 diode
R24282 N24281 N24282 10
D24282 N24282 0 diode
R24283 N24282 N24283 10
D24283 N24283 0 diode
R24284 N24283 N24284 10
D24284 N24284 0 diode
R24285 N24284 N24285 10
D24285 N24285 0 diode
R24286 N24285 N24286 10
D24286 N24286 0 diode
R24287 N24286 N24287 10
D24287 N24287 0 diode
R24288 N24287 N24288 10
D24288 N24288 0 diode
R24289 N24288 N24289 10
D24289 N24289 0 diode
R24290 N24289 N24290 10
D24290 N24290 0 diode
R24291 N24290 N24291 10
D24291 N24291 0 diode
R24292 N24291 N24292 10
D24292 N24292 0 diode
R24293 N24292 N24293 10
D24293 N24293 0 diode
R24294 N24293 N24294 10
D24294 N24294 0 diode
R24295 N24294 N24295 10
D24295 N24295 0 diode
R24296 N24295 N24296 10
D24296 N24296 0 diode
R24297 N24296 N24297 10
D24297 N24297 0 diode
R24298 N24297 N24298 10
D24298 N24298 0 diode
R24299 N24298 N24299 10
D24299 N24299 0 diode
R24300 N24299 N24300 10
D24300 N24300 0 diode
R24301 N24300 N24301 10
D24301 N24301 0 diode
R24302 N24301 N24302 10
D24302 N24302 0 diode
R24303 N24302 N24303 10
D24303 N24303 0 diode
R24304 N24303 N24304 10
D24304 N24304 0 diode
R24305 N24304 N24305 10
D24305 N24305 0 diode
R24306 N24305 N24306 10
D24306 N24306 0 diode
R24307 N24306 N24307 10
D24307 N24307 0 diode
R24308 N24307 N24308 10
D24308 N24308 0 diode
R24309 N24308 N24309 10
D24309 N24309 0 diode
R24310 N24309 N24310 10
D24310 N24310 0 diode
R24311 N24310 N24311 10
D24311 N24311 0 diode
R24312 N24311 N24312 10
D24312 N24312 0 diode
R24313 N24312 N24313 10
D24313 N24313 0 diode
R24314 N24313 N24314 10
D24314 N24314 0 diode
R24315 N24314 N24315 10
D24315 N24315 0 diode
R24316 N24315 N24316 10
D24316 N24316 0 diode
R24317 N24316 N24317 10
D24317 N24317 0 diode
R24318 N24317 N24318 10
D24318 N24318 0 diode
R24319 N24318 N24319 10
D24319 N24319 0 diode
R24320 N24319 N24320 10
D24320 N24320 0 diode
R24321 N24320 N24321 10
D24321 N24321 0 diode
R24322 N24321 N24322 10
D24322 N24322 0 diode
R24323 N24322 N24323 10
D24323 N24323 0 diode
R24324 N24323 N24324 10
D24324 N24324 0 diode
R24325 N24324 N24325 10
D24325 N24325 0 diode
R24326 N24325 N24326 10
D24326 N24326 0 diode
R24327 N24326 N24327 10
D24327 N24327 0 diode
R24328 N24327 N24328 10
D24328 N24328 0 diode
R24329 N24328 N24329 10
D24329 N24329 0 diode
R24330 N24329 N24330 10
D24330 N24330 0 diode
R24331 N24330 N24331 10
D24331 N24331 0 diode
R24332 N24331 N24332 10
D24332 N24332 0 diode
R24333 N24332 N24333 10
D24333 N24333 0 diode
R24334 N24333 N24334 10
D24334 N24334 0 diode
R24335 N24334 N24335 10
D24335 N24335 0 diode
R24336 N24335 N24336 10
D24336 N24336 0 diode
R24337 N24336 N24337 10
D24337 N24337 0 diode
R24338 N24337 N24338 10
D24338 N24338 0 diode
R24339 N24338 N24339 10
D24339 N24339 0 diode
R24340 N24339 N24340 10
D24340 N24340 0 diode
R24341 N24340 N24341 10
D24341 N24341 0 diode
R24342 N24341 N24342 10
D24342 N24342 0 diode
R24343 N24342 N24343 10
D24343 N24343 0 diode
R24344 N24343 N24344 10
D24344 N24344 0 diode
R24345 N24344 N24345 10
D24345 N24345 0 diode
R24346 N24345 N24346 10
D24346 N24346 0 diode
R24347 N24346 N24347 10
D24347 N24347 0 diode
R24348 N24347 N24348 10
D24348 N24348 0 diode
R24349 N24348 N24349 10
D24349 N24349 0 diode
R24350 N24349 N24350 10
D24350 N24350 0 diode
R24351 N24350 N24351 10
D24351 N24351 0 diode
R24352 N24351 N24352 10
D24352 N24352 0 diode
R24353 N24352 N24353 10
D24353 N24353 0 diode
R24354 N24353 N24354 10
D24354 N24354 0 diode
R24355 N24354 N24355 10
D24355 N24355 0 diode
R24356 N24355 N24356 10
D24356 N24356 0 diode
R24357 N24356 N24357 10
D24357 N24357 0 diode
R24358 N24357 N24358 10
D24358 N24358 0 diode
R24359 N24358 N24359 10
D24359 N24359 0 diode
R24360 N24359 N24360 10
D24360 N24360 0 diode
R24361 N24360 N24361 10
D24361 N24361 0 diode
R24362 N24361 N24362 10
D24362 N24362 0 diode
R24363 N24362 N24363 10
D24363 N24363 0 diode
R24364 N24363 N24364 10
D24364 N24364 0 diode
R24365 N24364 N24365 10
D24365 N24365 0 diode
R24366 N24365 N24366 10
D24366 N24366 0 diode
R24367 N24366 N24367 10
D24367 N24367 0 diode
R24368 N24367 N24368 10
D24368 N24368 0 diode
R24369 N24368 N24369 10
D24369 N24369 0 diode
R24370 N24369 N24370 10
D24370 N24370 0 diode
R24371 N24370 N24371 10
D24371 N24371 0 diode
R24372 N24371 N24372 10
D24372 N24372 0 diode
R24373 N24372 N24373 10
D24373 N24373 0 diode
R24374 N24373 N24374 10
D24374 N24374 0 diode
R24375 N24374 N24375 10
D24375 N24375 0 diode
R24376 N24375 N24376 10
D24376 N24376 0 diode
R24377 N24376 N24377 10
D24377 N24377 0 diode
R24378 N24377 N24378 10
D24378 N24378 0 diode
R24379 N24378 N24379 10
D24379 N24379 0 diode
R24380 N24379 N24380 10
D24380 N24380 0 diode
R24381 N24380 N24381 10
D24381 N24381 0 diode
R24382 N24381 N24382 10
D24382 N24382 0 diode
R24383 N24382 N24383 10
D24383 N24383 0 diode
R24384 N24383 N24384 10
D24384 N24384 0 diode
R24385 N24384 N24385 10
D24385 N24385 0 diode
R24386 N24385 N24386 10
D24386 N24386 0 diode
R24387 N24386 N24387 10
D24387 N24387 0 diode
R24388 N24387 N24388 10
D24388 N24388 0 diode
R24389 N24388 N24389 10
D24389 N24389 0 diode
R24390 N24389 N24390 10
D24390 N24390 0 diode
R24391 N24390 N24391 10
D24391 N24391 0 diode
R24392 N24391 N24392 10
D24392 N24392 0 diode
R24393 N24392 N24393 10
D24393 N24393 0 diode
R24394 N24393 N24394 10
D24394 N24394 0 diode
R24395 N24394 N24395 10
D24395 N24395 0 diode
R24396 N24395 N24396 10
D24396 N24396 0 diode
R24397 N24396 N24397 10
D24397 N24397 0 diode
R24398 N24397 N24398 10
D24398 N24398 0 diode
R24399 N24398 N24399 10
D24399 N24399 0 diode
R24400 N24399 N24400 10
D24400 N24400 0 diode
R24401 N24400 N24401 10
D24401 N24401 0 diode
R24402 N24401 N24402 10
D24402 N24402 0 diode
R24403 N24402 N24403 10
D24403 N24403 0 diode
R24404 N24403 N24404 10
D24404 N24404 0 diode
R24405 N24404 N24405 10
D24405 N24405 0 diode
R24406 N24405 N24406 10
D24406 N24406 0 diode
R24407 N24406 N24407 10
D24407 N24407 0 diode
R24408 N24407 N24408 10
D24408 N24408 0 diode
R24409 N24408 N24409 10
D24409 N24409 0 diode
R24410 N24409 N24410 10
D24410 N24410 0 diode
R24411 N24410 N24411 10
D24411 N24411 0 diode
R24412 N24411 N24412 10
D24412 N24412 0 diode
R24413 N24412 N24413 10
D24413 N24413 0 diode
R24414 N24413 N24414 10
D24414 N24414 0 diode
R24415 N24414 N24415 10
D24415 N24415 0 diode
R24416 N24415 N24416 10
D24416 N24416 0 diode
R24417 N24416 N24417 10
D24417 N24417 0 diode
R24418 N24417 N24418 10
D24418 N24418 0 diode
R24419 N24418 N24419 10
D24419 N24419 0 diode
R24420 N24419 N24420 10
D24420 N24420 0 diode
R24421 N24420 N24421 10
D24421 N24421 0 diode
R24422 N24421 N24422 10
D24422 N24422 0 diode
R24423 N24422 N24423 10
D24423 N24423 0 diode
R24424 N24423 N24424 10
D24424 N24424 0 diode
R24425 N24424 N24425 10
D24425 N24425 0 diode
R24426 N24425 N24426 10
D24426 N24426 0 diode
R24427 N24426 N24427 10
D24427 N24427 0 diode
R24428 N24427 N24428 10
D24428 N24428 0 diode
R24429 N24428 N24429 10
D24429 N24429 0 diode
R24430 N24429 N24430 10
D24430 N24430 0 diode
R24431 N24430 N24431 10
D24431 N24431 0 diode
R24432 N24431 N24432 10
D24432 N24432 0 diode
R24433 N24432 N24433 10
D24433 N24433 0 diode
R24434 N24433 N24434 10
D24434 N24434 0 diode
R24435 N24434 N24435 10
D24435 N24435 0 diode
R24436 N24435 N24436 10
D24436 N24436 0 diode
R24437 N24436 N24437 10
D24437 N24437 0 diode
R24438 N24437 N24438 10
D24438 N24438 0 diode
R24439 N24438 N24439 10
D24439 N24439 0 diode
R24440 N24439 N24440 10
D24440 N24440 0 diode
R24441 N24440 N24441 10
D24441 N24441 0 diode
R24442 N24441 N24442 10
D24442 N24442 0 diode
R24443 N24442 N24443 10
D24443 N24443 0 diode
R24444 N24443 N24444 10
D24444 N24444 0 diode
R24445 N24444 N24445 10
D24445 N24445 0 diode
R24446 N24445 N24446 10
D24446 N24446 0 diode
R24447 N24446 N24447 10
D24447 N24447 0 diode
R24448 N24447 N24448 10
D24448 N24448 0 diode
R24449 N24448 N24449 10
D24449 N24449 0 diode
R24450 N24449 N24450 10
D24450 N24450 0 diode
R24451 N24450 N24451 10
D24451 N24451 0 diode
R24452 N24451 N24452 10
D24452 N24452 0 diode
R24453 N24452 N24453 10
D24453 N24453 0 diode
R24454 N24453 N24454 10
D24454 N24454 0 diode
R24455 N24454 N24455 10
D24455 N24455 0 diode
R24456 N24455 N24456 10
D24456 N24456 0 diode
R24457 N24456 N24457 10
D24457 N24457 0 diode
R24458 N24457 N24458 10
D24458 N24458 0 diode
R24459 N24458 N24459 10
D24459 N24459 0 diode
R24460 N24459 N24460 10
D24460 N24460 0 diode
R24461 N24460 N24461 10
D24461 N24461 0 diode
R24462 N24461 N24462 10
D24462 N24462 0 diode
R24463 N24462 N24463 10
D24463 N24463 0 diode
R24464 N24463 N24464 10
D24464 N24464 0 diode
R24465 N24464 N24465 10
D24465 N24465 0 diode
R24466 N24465 N24466 10
D24466 N24466 0 diode
R24467 N24466 N24467 10
D24467 N24467 0 diode
R24468 N24467 N24468 10
D24468 N24468 0 diode
R24469 N24468 N24469 10
D24469 N24469 0 diode
R24470 N24469 N24470 10
D24470 N24470 0 diode
R24471 N24470 N24471 10
D24471 N24471 0 diode
R24472 N24471 N24472 10
D24472 N24472 0 diode
R24473 N24472 N24473 10
D24473 N24473 0 diode
R24474 N24473 N24474 10
D24474 N24474 0 diode
R24475 N24474 N24475 10
D24475 N24475 0 diode
R24476 N24475 N24476 10
D24476 N24476 0 diode
R24477 N24476 N24477 10
D24477 N24477 0 diode
R24478 N24477 N24478 10
D24478 N24478 0 diode
R24479 N24478 N24479 10
D24479 N24479 0 diode
R24480 N24479 N24480 10
D24480 N24480 0 diode
R24481 N24480 N24481 10
D24481 N24481 0 diode
R24482 N24481 N24482 10
D24482 N24482 0 diode
R24483 N24482 N24483 10
D24483 N24483 0 diode
R24484 N24483 N24484 10
D24484 N24484 0 diode
R24485 N24484 N24485 10
D24485 N24485 0 diode
R24486 N24485 N24486 10
D24486 N24486 0 diode
R24487 N24486 N24487 10
D24487 N24487 0 diode
R24488 N24487 N24488 10
D24488 N24488 0 diode
R24489 N24488 N24489 10
D24489 N24489 0 diode
R24490 N24489 N24490 10
D24490 N24490 0 diode
R24491 N24490 N24491 10
D24491 N24491 0 diode
R24492 N24491 N24492 10
D24492 N24492 0 diode
R24493 N24492 N24493 10
D24493 N24493 0 diode
R24494 N24493 N24494 10
D24494 N24494 0 diode
R24495 N24494 N24495 10
D24495 N24495 0 diode
R24496 N24495 N24496 10
D24496 N24496 0 diode
R24497 N24496 N24497 10
D24497 N24497 0 diode
R24498 N24497 N24498 10
D24498 N24498 0 diode
R24499 N24498 N24499 10
D24499 N24499 0 diode
R24500 N24499 N24500 10
D24500 N24500 0 diode
R24501 N24500 N24501 10
D24501 N24501 0 diode
R24502 N24501 N24502 10
D24502 N24502 0 diode
R24503 N24502 N24503 10
D24503 N24503 0 diode
R24504 N24503 N24504 10
D24504 N24504 0 diode
R24505 N24504 N24505 10
D24505 N24505 0 diode
R24506 N24505 N24506 10
D24506 N24506 0 diode
R24507 N24506 N24507 10
D24507 N24507 0 diode
R24508 N24507 N24508 10
D24508 N24508 0 diode
R24509 N24508 N24509 10
D24509 N24509 0 diode
R24510 N24509 N24510 10
D24510 N24510 0 diode
R24511 N24510 N24511 10
D24511 N24511 0 diode
R24512 N24511 N24512 10
D24512 N24512 0 diode
R24513 N24512 N24513 10
D24513 N24513 0 diode
R24514 N24513 N24514 10
D24514 N24514 0 diode
R24515 N24514 N24515 10
D24515 N24515 0 diode
R24516 N24515 N24516 10
D24516 N24516 0 diode
R24517 N24516 N24517 10
D24517 N24517 0 diode
R24518 N24517 N24518 10
D24518 N24518 0 diode
R24519 N24518 N24519 10
D24519 N24519 0 diode
R24520 N24519 N24520 10
D24520 N24520 0 diode
R24521 N24520 N24521 10
D24521 N24521 0 diode
R24522 N24521 N24522 10
D24522 N24522 0 diode
R24523 N24522 N24523 10
D24523 N24523 0 diode
R24524 N24523 N24524 10
D24524 N24524 0 diode
R24525 N24524 N24525 10
D24525 N24525 0 diode
R24526 N24525 N24526 10
D24526 N24526 0 diode
R24527 N24526 N24527 10
D24527 N24527 0 diode
R24528 N24527 N24528 10
D24528 N24528 0 diode
R24529 N24528 N24529 10
D24529 N24529 0 diode
R24530 N24529 N24530 10
D24530 N24530 0 diode
R24531 N24530 N24531 10
D24531 N24531 0 diode
R24532 N24531 N24532 10
D24532 N24532 0 diode
R24533 N24532 N24533 10
D24533 N24533 0 diode
R24534 N24533 N24534 10
D24534 N24534 0 diode
R24535 N24534 N24535 10
D24535 N24535 0 diode
R24536 N24535 N24536 10
D24536 N24536 0 diode
R24537 N24536 N24537 10
D24537 N24537 0 diode
R24538 N24537 N24538 10
D24538 N24538 0 diode
R24539 N24538 N24539 10
D24539 N24539 0 diode
R24540 N24539 N24540 10
D24540 N24540 0 diode
R24541 N24540 N24541 10
D24541 N24541 0 diode
R24542 N24541 N24542 10
D24542 N24542 0 diode
R24543 N24542 N24543 10
D24543 N24543 0 diode
R24544 N24543 N24544 10
D24544 N24544 0 diode
R24545 N24544 N24545 10
D24545 N24545 0 diode
R24546 N24545 N24546 10
D24546 N24546 0 diode
R24547 N24546 N24547 10
D24547 N24547 0 diode
R24548 N24547 N24548 10
D24548 N24548 0 diode
R24549 N24548 N24549 10
D24549 N24549 0 diode
R24550 N24549 N24550 10
D24550 N24550 0 diode
R24551 N24550 N24551 10
D24551 N24551 0 diode
R24552 N24551 N24552 10
D24552 N24552 0 diode
R24553 N24552 N24553 10
D24553 N24553 0 diode
R24554 N24553 N24554 10
D24554 N24554 0 diode
R24555 N24554 N24555 10
D24555 N24555 0 diode
R24556 N24555 N24556 10
D24556 N24556 0 diode
R24557 N24556 N24557 10
D24557 N24557 0 diode
R24558 N24557 N24558 10
D24558 N24558 0 diode
R24559 N24558 N24559 10
D24559 N24559 0 diode
R24560 N24559 N24560 10
D24560 N24560 0 diode
R24561 N24560 N24561 10
D24561 N24561 0 diode
R24562 N24561 N24562 10
D24562 N24562 0 diode
R24563 N24562 N24563 10
D24563 N24563 0 diode
R24564 N24563 N24564 10
D24564 N24564 0 diode
R24565 N24564 N24565 10
D24565 N24565 0 diode
R24566 N24565 N24566 10
D24566 N24566 0 diode
R24567 N24566 N24567 10
D24567 N24567 0 diode
R24568 N24567 N24568 10
D24568 N24568 0 diode
R24569 N24568 N24569 10
D24569 N24569 0 diode
R24570 N24569 N24570 10
D24570 N24570 0 diode
R24571 N24570 N24571 10
D24571 N24571 0 diode
R24572 N24571 N24572 10
D24572 N24572 0 diode
R24573 N24572 N24573 10
D24573 N24573 0 diode
R24574 N24573 N24574 10
D24574 N24574 0 diode
R24575 N24574 N24575 10
D24575 N24575 0 diode
R24576 N24575 N24576 10
D24576 N24576 0 diode
R24577 N24576 N24577 10
D24577 N24577 0 diode
R24578 N24577 N24578 10
D24578 N24578 0 diode
R24579 N24578 N24579 10
D24579 N24579 0 diode
R24580 N24579 N24580 10
D24580 N24580 0 diode
R24581 N24580 N24581 10
D24581 N24581 0 diode
R24582 N24581 N24582 10
D24582 N24582 0 diode
R24583 N24582 N24583 10
D24583 N24583 0 diode
R24584 N24583 N24584 10
D24584 N24584 0 diode
R24585 N24584 N24585 10
D24585 N24585 0 diode
R24586 N24585 N24586 10
D24586 N24586 0 diode
R24587 N24586 N24587 10
D24587 N24587 0 diode
R24588 N24587 N24588 10
D24588 N24588 0 diode
R24589 N24588 N24589 10
D24589 N24589 0 diode
R24590 N24589 N24590 10
D24590 N24590 0 diode
R24591 N24590 N24591 10
D24591 N24591 0 diode
R24592 N24591 N24592 10
D24592 N24592 0 diode
R24593 N24592 N24593 10
D24593 N24593 0 diode
R24594 N24593 N24594 10
D24594 N24594 0 diode
R24595 N24594 N24595 10
D24595 N24595 0 diode
R24596 N24595 N24596 10
D24596 N24596 0 diode
R24597 N24596 N24597 10
D24597 N24597 0 diode
R24598 N24597 N24598 10
D24598 N24598 0 diode
R24599 N24598 N24599 10
D24599 N24599 0 diode
R24600 N24599 N24600 10
D24600 N24600 0 diode
R24601 N24600 N24601 10
D24601 N24601 0 diode
R24602 N24601 N24602 10
D24602 N24602 0 diode
R24603 N24602 N24603 10
D24603 N24603 0 diode
R24604 N24603 N24604 10
D24604 N24604 0 diode
R24605 N24604 N24605 10
D24605 N24605 0 diode
R24606 N24605 N24606 10
D24606 N24606 0 diode
R24607 N24606 N24607 10
D24607 N24607 0 diode
R24608 N24607 N24608 10
D24608 N24608 0 diode
R24609 N24608 N24609 10
D24609 N24609 0 diode
R24610 N24609 N24610 10
D24610 N24610 0 diode
R24611 N24610 N24611 10
D24611 N24611 0 diode
R24612 N24611 N24612 10
D24612 N24612 0 diode
R24613 N24612 N24613 10
D24613 N24613 0 diode
R24614 N24613 N24614 10
D24614 N24614 0 diode
R24615 N24614 N24615 10
D24615 N24615 0 diode
R24616 N24615 N24616 10
D24616 N24616 0 diode
R24617 N24616 N24617 10
D24617 N24617 0 diode
R24618 N24617 N24618 10
D24618 N24618 0 diode
R24619 N24618 N24619 10
D24619 N24619 0 diode
R24620 N24619 N24620 10
D24620 N24620 0 diode
R24621 N24620 N24621 10
D24621 N24621 0 diode
R24622 N24621 N24622 10
D24622 N24622 0 diode
R24623 N24622 N24623 10
D24623 N24623 0 diode
R24624 N24623 N24624 10
D24624 N24624 0 diode
R24625 N24624 N24625 10
D24625 N24625 0 diode
R24626 N24625 N24626 10
D24626 N24626 0 diode
R24627 N24626 N24627 10
D24627 N24627 0 diode
R24628 N24627 N24628 10
D24628 N24628 0 diode
R24629 N24628 N24629 10
D24629 N24629 0 diode
R24630 N24629 N24630 10
D24630 N24630 0 diode
R24631 N24630 N24631 10
D24631 N24631 0 diode
R24632 N24631 N24632 10
D24632 N24632 0 diode
R24633 N24632 N24633 10
D24633 N24633 0 diode
R24634 N24633 N24634 10
D24634 N24634 0 diode
R24635 N24634 N24635 10
D24635 N24635 0 diode
R24636 N24635 N24636 10
D24636 N24636 0 diode
R24637 N24636 N24637 10
D24637 N24637 0 diode
R24638 N24637 N24638 10
D24638 N24638 0 diode
R24639 N24638 N24639 10
D24639 N24639 0 diode
R24640 N24639 N24640 10
D24640 N24640 0 diode
R24641 N24640 N24641 10
D24641 N24641 0 diode
R24642 N24641 N24642 10
D24642 N24642 0 diode
R24643 N24642 N24643 10
D24643 N24643 0 diode
R24644 N24643 N24644 10
D24644 N24644 0 diode
R24645 N24644 N24645 10
D24645 N24645 0 diode
R24646 N24645 N24646 10
D24646 N24646 0 diode
R24647 N24646 N24647 10
D24647 N24647 0 diode
R24648 N24647 N24648 10
D24648 N24648 0 diode
R24649 N24648 N24649 10
D24649 N24649 0 diode
R24650 N24649 N24650 10
D24650 N24650 0 diode
R24651 N24650 N24651 10
D24651 N24651 0 diode
R24652 N24651 N24652 10
D24652 N24652 0 diode
R24653 N24652 N24653 10
D24653 N24653 0 diode
R24654 N24653 N24654 10
D24654 N24654 0 diode
R24655 N24654 N24655 10
D24655 N24655 0 diode
R24656 N24655 N24656 10
D24656 N24656 0 diode
R24657 N24656 N24657 10
D24657 N24657 0 diode
R24658 N24657 N24658 10
D24658 N24658 0 diode
R24659 N24658 N24659 10
D24659 N24659 0 diode
R24660 N24659 N24660 10
D24660 N24660 0 diode
R24661 N24660 N24661 10
D24661 N24661 0 diode
R24662 N24661 N24662 10
D24662 N24662 0 diode
R24663 N24662 N24663 10
D24663 N24663 0 diode
R24664 N24663 N24664 10
D24664 N24664 0 diode
R24665 N24664 N24665 10
D24665 N24665 0 diode
R24666 N24665 N24666 10
D24666 N24666 0 diode
R24667 N24666 N24667 10
D24667 N24667 0 diode
R24668 N24667 N24668 10
D24668 N24668 0 diode
R24669 N24668 N24669 10
D24669 N24669 0 diode
R24670 N24669 N24670 10
D24670 N24670 0 diode
R24671 N24670 N24671 10
D24671 N24671 0 diode
R24672 N24671 N24672 10
D24672 N24672 0 diode
R24673 N24672 N24673 10
D24673 N24673 0 diode
R24674 N24673 N24674 10
D24674 N24674 0 diode
R24675 N24674 N24675 10
D24675 N24675 0 diode
R24676 N24675 N24676 10
D24676 N24676 0 diode
R24677 N24676 N24677 10
D24677 N24677 0 diode
R24678 N24677 N24678 10
D24678 N24678 0 diode
R24679 N24678 N24679 10
D24679 N24679 0 diode
R24680 N24679 N24680 10
D24680 N24680 0 diode
R24681 N24680 N24681 10
D24681 N24681 0 diode
R24682 N24681 N24682 10
D24682 N24682 0 diode
R24683 N24682 N24683 10
D24683 N24683 0 diode
R24684 N24683 N24684 10
D24684 N24684 0 diode
R24685 N24684 N24685 10
D24685 N24685 0 diode
R24686 N24685 N24686 10
D24686 N24686 0 diode
R24687 N24686 N24687 10
D24687 N24687 0 diode
R24688 N24687 N24688 10
D24688 N24688 0 diode
R24689 N24688 N24689 10
D24689 N24689 0 diode
R24690 N24689 N24690 10
D24690 N24690 0 diode
R24691 N24690 N24691 10
D24691 N24691 0 diode
R24692 N24691 N24692 10
D24692 N24692 0 diode
R24693 N24692 N24693 10
D24693 N24693 0 diode
R24694 N24693 N24694 10
D24694 N24694 0 diode
R24695 N24694 N24695 10
D24695 N24695 0 diode
R24696 N24695 N24696 10
D24696 N24696 0 diode
R24697 N24696 N24697 10
D24697 N24697 0 diode
R24698 N24697 N24698 10
D24698 N24698 0 diode
R24699 N24698 N24699 10
D24699 N24699 0 diode
R24700 N24699 N24700 10
D24700 N24700 0 diode
R24701 N24700 N24701 10
D24701 N24701 0 diode
R24702 N24701 N24702 10
D24702 N24702 0 diode
R24703 N24702 N24703 10
D24703 N24703 0 diode
R24704 N24703 N24704 10
D24704 N24704 0 diode
R24705 N24704 N24705 10
D24705 N24705 0 diode
R24706 N24705 N24706 10
D24706 N24706 0 diode
R24707 N24706 N24707 10
D24707 N24707 0 diode
R24708 N24707 N24708 10
D24708 N24708 0 diode
R24709 N24708 N24709 10
D24709 N24709 0 diode
R24710 N24709 N24710 10
D24710 N24710 0 diode
R24711 N24710 N24711 10
D24711 N24711 0 diode
R24712 N24711 N24712 10
D24712 N24712 0 diode
R24713 N24712 N24713 10
D24713 N24713 0 diode
R24714 N24713 N24714 10
D24714 N24714 0 diode
R24715 N24714 N24715 10
D24715 N24715 0 diode
R24716 N24715 N24716 10
D24716 N24716 0 diode
R24717 N24716 N24717 10
D24717 N24717 0 diode
R24718 N24717 N24718 10
D24718 N24718 0 diode
R24719 N24718 N24719 10
D24719 N24719 0 diode
R24720 N24719 N24720 10
D24720 N24720 0 diode
R24721 N24720 N24721 10
D24721 N24721 0 diode
R24722 N24721 N24722 10
D24722 N24722 0 diode
R24723 N24722 N24723 10
D24723 N24723 0 diode
R24724 N24723 N24724 10
D24724 N24724 0 diode
R24725 N24724 N24725 10
D24725 N24725 0 diode
R24726 N24725 N24726 10
D24726 N24726 0 diode
R24727 N24726 N24727 10
D24727 N24727 0 diode
R24728 N24727 N24728 10
D24728 N24728 0 diode
R24729 N24728 N24729 10
D24729 N24729 0 diode
R24730 N24729 N24730 10
D24730 N24730 0 diode
R24731 N24730 N24731 10
D24731 N24731 0 diode
R24732 N24731 N24732 10
D24732 N24732 0 diode
R24733 N24732 N24733 10
D24733 N24733 0 diode
R24734 N24733 N24734 10
D24734 N24734 0 diode
R24735 N24734 N24735 10
D24735 N24735 0 diode
R24736 N24735 N24736 10
D24736 N24736 0 diode
R24737 N24736 N24737 10
D24737 N24737 0 diode
R24738 N24737 N24738 10
D24738 N24738 0 diode
R24739 N24738 N24739 10
D24739 N24739 0 diode
R24740 N24739 N24740 10
D24740 N24740 0 diode
R24741 N24740 N24741 10
D24741 N24741 0 diode
R24742 N24741 N24742 10
D24742 N24742 0 diode
R24743 N24742 N24743 10
D24743 N24743 0 diode
R24744 N24743 N24744 10
D24744 N24744 0 diode
R24745 N24744 N24745 10
D24745 N24745 0 diode
R24746 N24745 N24746 10
D24746 N24746 0 diode
R24747 N24746 N24747 10
D24747 N24747 0 diode
R24748 N24747 N24748 10
D24748 N24748 0 diode
R24749 N24748 N24749 10
D24749 N24749 0 diode
R24750 N24749 N24750 10
D24750 N24750 0 diode
R24751 N24750 N24751 10
D24751 N24751 0 diode
R24752 N24751 N24752 10
D24752 N24752 0 diode
R24753 N24752 N24753 10
D24753 N24753 0 diode
R24754 N24753 N24754 10
D24754 N24754 0 diode
R24755 N24754 N24755 10
D24755 N24755 0 diode
R24756 N24755 N24756 10
D24756 N24756 0 diode
R24757 N24756 N24757 10
D24757 N24757 0 diode
R24758 N24757 N24758 10
D24758 N24758 0 diode
R24759 N24758 N24759 10
D24759 N24759 0 diode
R24760 N24759 N24760 10
D24760 N24760 0 diode
R24761 N24760 N24761 10
D24761 N24761 0 diode
R24762 N24761 N24762 10
D24762 N24762 0 diode
R24763 N24762 N24763 10
D24763 N24763 0 diode
R24764 N24763 N24764 10
D24764 N24764 0 diode
R24765 N24764 N24765 10
D24765 N24765 0 diode
R24766 N24765 N24766 10
D24766 N24766 0 diode
R24767 N24766 N24767 10
D24767 N24767 0 diode
R24768 N24767 N24768 10
D24768 N24768 0 diode
R24769 N24768 N24769 10
D24769 N24769 0 diode
R24770 N24769 N24770 10
D24770 N24770 0 diode
R24771 N24770 N24771 10
D24771 N24771 0 diode
R24772 N24771 N24772 10
D24772 N24772 0 diode
R24773 N24772 N24773 10
D24773 N24773 0 diode
R24774 N24773 N24774 10
D24774 N24774 0 diode
R24775 N24774 N24775 10
D24775 N24775 0 diode
R24776 N24775 N24776 10
D24776 N24776 0 diode
R24777 N24776 N24777 10
D24777 N24777 0 diode
R24778 N24777 N24778 10
D24778 N24778 0 diode
R24779 N24778 N24779 10
D24779 N24779 0 diode
R24780 N24779 N24780 10
D24780 N24780 0 diode
R24781 N24780 N24781 10
D24781 N24781 0 diode
R24782 N24781 N24782 10
D24782 N24782 0 diode
R24783 N24782 N24783 10
D24783 N24783 0 diode
R24784 N24783 N24784 10
D24784 N24784 0 diode
R24785 N24784 N24785 10
D24785 N24785 0 diode
R24786 N24785 N24786 10
D24786 N24786 0 diode
R24787 N24786 N24787 10
D24787 N24787 0 diode
R24788 N24787 N24788 10
D24788 N24788 0 diode
R24789 N24788 N24789 10
D24789 N24789 0 diode
R24790 N24789 N24790 10
D24790 N24790 0 diode
R24791 N24790 N24791 10
D24791 N24791 0 diode
R24792 N24791 N24792 10
D24792 N24792 0 diode
R24793 N24792 N24793 10
D24793 N24793 0 diode
R24794 N24793 N24794 10
D24794 N24794 0 diode
R24795 N24794 N24795 10
D24795 N24795 0 diode
R24796 N24795 N24796 10
D24796 N24796 0 diode
R24797 N24796 N24797 10
D24797 N24797 0 diode
R24798 N24797 N24798 10
D24798 N24798 0 diode
R24799 N24798 N24799 10
D24799 N24799 0 diode
R24800 N24799 N24800 10
D24800 N24800 0 diode
R24801 N24800 N24801 10
D24801 N24801 0 diode
R24802 N24801 N24802 10
D24802 N24802 0 diode
R24803 N24802 N24803 10
D24803 N24803 0 diode
R24804 N24803 N24804 10
D24804 N24804 0 diode
R24805 N24804 N24805 10
D24805 N24805 0 diode
R24806 N24805 N24806 10
D24806 N24806 0 diode
R24807 N24806 N24807 10
D24807 N24807 0 diode
R24808 N24807 N24808 10
D24808 N24808 0 diode
R24809 N24808 N24809 10
D24809 N24809 0 diode
R24810 N24809 N24810 10
D24810 N24810 0 diode
R24811 N24810 N24811 10
D24811 N24811 0 diode
R24812 N24811 N24812 10
D24812 N24812 0 diode
R24813 N24812 N24813 10
D24813 N24813 0 diode
R24814 N24813 N24814 10
D24814 N24814 0 diode
R24815 N24814 N24815 10
D24815 N24815 0 diode
R24816 N24815 N24816 10
D24816 N24816 0 diode
R24817 N24816 N24817 10
D24817 N24817 0 diode
R24818 N24817 N24818 10
D24818 N24818 0 diode
R24819 N24818 N24819 10
D24819 N24819 0 diode
R24820 N24819 N24820 10
D24820 N24820 0 diode
R24821 N24820 N24821 10
D24821 N24821 0 diode
R24822 N24821 N24822 10
D24822 N24822 0 diode
R24823 N24822 N24823 10
D24823 N24823 0 diode
R24824 N24823 N24824 10
D24824 N24824 0 diode
R24825 N24824 N24825 10
D24825 N24825 0 diode
R24826 N24825 N24826 10
D24826 N24826 0 diode
R24827 N24826 N24827 10
D24827 N24827 0 diode
R24828 N24827 N24828 10
D24828 N24828 0 diode
R24829 N24828 N24829 10
D24829 N24829 0 diode
R24830 N24829 N24830 10
D24830 N24830 0 diode
R24831 N24830 N24831 10
D24831 N24831 0 diode
R24832 N24831 N24832 10
D24832 N24832 0 diode
R24833 N24832 N24833 10
D24833 N24833 0 diode
R24834 N24833 N24834 10
D24834 N24834 0 diode
R24835 N24834 N24835 10
D24835 N24835 0 diode
R24836 N24835 N24836 10
D24836 N24836 0 diode
R24837 N24836 N24837 10
D24837 N24837 0 diode
R24838 N24837 N24838 10
D24838 N24838 0 diode
R24839 N24838 N24839 10
D24839 N24839 0 diode
R24840 N24839 N24840 10
D24840 N24840 0 diode
R24841 N24840 N24841 10
D24841 N24841 0 diode
R24842 N24841 N24842 10
D24842 N24842 0 diode
R24843 N24842 N24843 10
D24843 N24843 0 diode
R24844 N24843 N24844 10
D24844 N24844 0 diode
R24845 N24844 N24845 10
D24845 N24845 0 diode
R24846 N24845 N24846 10
D24846 N24846 0 diode
R24847 N24846 N24847 10
D24847 N24847 0 diode
R24848 N24847 N24848 10
D24848 N24848 0 diode
R24849 N24848 N24849 10
D24849 N24849 0 diode
R24850 N24849 N24850 10
D24850 N24850 0 diode
R24851 N24850 N24851 10
D24851 N24851 0 diode
R24852 N24851 N24852 10
D24852 N24852 0 diode
R24853 N24852 N24853 10
D24853 N24853 0 diode
R24854 N24853 N24854 10
D24854 N24854 0 diode
R24855 N24854 N24855 10
D24855 N24855 0 diode
R24856 N24855 N24856 10
D24856 N24856 0 diode
R24857 N24856 N24857 10
D24857 N24857 0 diode
R24858 N24857 N24858 10
D24858 N24858 0 diode
R24859 N24858 N24859 10
D24859 N24859 0 diode
R24860 N24859 N24860 10
D24860 N24860 0 diode
R24861 N24860 N24861 10
D24861 N24861 0 diode
R24862 N24861 N24862 10
D24862 N24862 0 diode
R24863 N24862 N24863 10
D24863 N24863 0 diode
R24864 N24863 N24864 10
D24864 N24864 0 diode
R24865 N24864 N24865 10
D24865 N24865 0 diode
R24866 N24865 N24866 10
D24866 N24866 0 diode
R24867 N24866 N24867 10
D24867 N24867 0 diode
R24868 N24867 N24868 10
D24868 N24868 0 diode
R24869 N24868 N24869 10
D24869 N24869 0 diode
R24870 N24869 N24870 10
D24870 N24870 0 diode
R24871 N24870 N24871 10
D24871 N24871 0 diode
R24872 N24871 N24872 10
D24872 N24872 0 diode
R24873 N24872 N24873 10
D24873 N24873 0 diode
R24874 N24873 N24874 10
D24874 N24874 0 diode
R24875 N24874 N24875 10
D24875 N24875 0 diode
R24876 N24875 N24876 10
D24876 N24876 0 diode
R24877 N24876 N24877 10
D24877 N24877 0 diode
R24878 N24877 N24878 10
D24878 N24878 0 diode
R24879 N24878 N24879 10
D24879 N24879 0 diode
R24880 N24879 N24880 10
D24880 N24880 0 diode
R24881 N24880 N24881 10
D24881 N24881 0 diode
R24882 N24881 N24882 10
D24882 N24882 0 diode
R24883 N24882 N24883 10
D24883 N24883 0 diode
R24884 N24883 N24884 10
D24884 N24884 0 diode
R24885 N24884 N24885 10
D24885 N24885 0 diode
R24886 N24885 N24886 10
D24886 N24886 0 diode
R24887 N24886 N24887 10
D24887 N24887 0 diode
R24888 N24887 N24888 10
D24888 N24888 0 diode
R24889 N24888 N24889 10
D24889 N24889 0 diode
R24890 N24889 N24890 10
D24890 N24890 0 diode
R24891 N24890 N24891 10
D24891 N24891 0 diode
R24892 N24891 N24892 10
D24892 N24892 0 diode
R24893 N24892 N24893 10
D24893 N24893 0 diode
R24894 N24893 N24894 10
D24894 N24894 0 diode
R24895 N24894 N24895 10
D24895 N24895 0 diode
R24896 N24895 N24896 10
D24896 N24896 0 diode
R24897 N24896 N24897 10
D24897 N24897 0 diode
R24898 N24897 N24898 10
D24898 N24898 0 diode
R24899 N24898 N24899 10
D24899 N24899 0 diode
R24900 N24899 N24900 10
D24900 N24900 0 diode
R24901 N24900 N24901 10
D24901 N24901 0 diode
R24902 N24901 N24902 10
D24902 N24902 0 diode
R24903 N24902 N24903 10
D24903 N24903 0 diode
R24904 N24903 N24904 10
D24904 N24904 0 diode
R24905 N24904 N24905 10
D24905 N24905 0 diode
R24906 N24905 N24906 10
D24906 N24906 0 diode
R24907 N24906 N24907 10
D24907 N24907 0 diode
R24908 N24907 N24908 10
D24908 N24908 0 diode
R24909 N24908 N24909 10
D24909 N24909 0 diode
R24910 N24909 N24910 10
D24910 N24910 0 diode
R24911 N24910 N24911 10
D24911 N24911 0 diode
R24912 N24911 N24912 10
D24912 N24912 0 diode
R24913 N24912 N24913 10
D24913 N24913 0 diode
R24914 N24913 N24914 10
D24914 N24914 0 diode
R24915 N24914 N24915 10
D24915 N24915 0 diode
R24916 N24915 N24916 10
D24916 N24916 0 diode
R24917 N24916 N24917 10
D24917 N24917 0 diode
R24918 N24917 N24918 10
D24918 N24918 0 diode
R24919 N24918 N24919 10
D24919 N24919 0 diode
R24920 N24919 N24920 10
D24920 N24920 0 diode
R24921 N24920 N24921 10
D24921 N24921 0 diode
R24922 N24921 N24922 10
D24922 N24922 0 diode
R24923 N24922 N24923 10
D24923 N24923 0 diode
R24924 N24923 N24924 10
D24924 N24924 0 diode
R24925 N24924 N24925 10
D24925 N24925 0 diode
R24926 N24925 N24926 10
D24926 N24926 0 diode
R24927 N24926 N24927 10
D24927 N24927 0 diode
R24928 N24927 N24928 10
D24928 N24928 0 diode
R24929 N24928 N24929 10
D24929 N24929 0 diode
R24930 N24929 N24930 10
D24930 N24930 0 diode
R24931 N24930 N24931 10
D24931 N24931 0 diode
R24932 N24931 N24932 10
D24932 N24932 0 diode
R24933 N24932 N24933 10
D24933 N24933 0 diode
R24934 N24933 N24934 10
D24934 N24934 0 diode
R24935 N24934 N24935 10
D24935 N24935 0 diode
R24936 N24935 N24936 10
D24936 N24936 0 diode
R24937 N24936 N24937 10
D24937 N24937 0 diode
R24938 N24937 N24938 10
D24938 N24938 0 diode
R24939 N24938 N24939 10
D24939 N24939 0 diode
R24940 N24939 N24940 10
D24940 N24940 0 diode
R24941 N24940 N24941 10
D24941 N24941 0 diode
R24942 N24941 N24942 10
D24942 N24942 0 diode
R24943 N24942 N24943 10
D24943 N24943 0 diode
R24944 N24943 N24944 10
D24944 N24944 0 diode
R24945 N24944 N24945 10
D24945 N24945 0 diode
R24946 N24945 N24946 10
D24946 N24946 0 diode
R24947 N24946 N24947 10
D24947 N24947 0 diode
R24948 N24947 N24948 10
D24948 N24948 0 diode
R24949 N24948 N24949 10
D24949 N24949 0 diode
R24950 N24949 N24950 10
D24950 N24950 0 diode
R24951 N24950 N24951 10
D24951 N24951 0 diode
R24952 N24951 N24952 10
D24952 N24952 0 diode
R24953 N24952 N24953 10
D24953 N24953 0 diode
R24954 N24953 N24954 10
D24954 N24954 0 diode
R24955 N24954 N24955 10
D24955 N24955 0 diode
R24956 N24955 N24956 10
D24956 N24956 0 diode
R24957 N24956 N24957 10
D24957 N24957 0 diode
R24958 N24957 N24958 10
D24958 N24958 0 diode
R24959 N24958 N24959 10
D24959 N24959 0 diode
R24960 N24959 N24960 10
D24960 N24960 0 diode
R24961 N24960 N24961 10
D24961 N24961 0 diode
R24962 N24961 N24962 10
D24962 N24962 0 diode
R24963 N24962 N24963 10
D24963 N24963 0 diode
R24964 N24963 N24964 10
D24964 N24964 0 diode
R24965 N24964 N24965 10
D24965 N24965 0 diode
R24966 N24965 N24966 10
D24966 N24966 0 diode
R24967 N24966 N24967 10
D24967 N24967 0 diode
R24968 N24967 N24968 10
D24968 N24968 0 diode
R24969 N24968 N24969 10
D24969 N24969 0 diode
R24970 N24969 N24970 10
D24970 N24970 0 diode
R24971 N24970 N24971 10
D24971 N24971 0 diode
R24972 N24971 N24972 10
D24972 N24972 0 diode
R24973 N24972 N24973 10
D24973 N24973 0 diode
R24974 N24973 N24974 10
D24974 N24974 0 diode
R24975 N24974 N24975 10
D24975 N24975 0 diode
R24976 N24975 N24976 10
D24976 N24976 0 diode
R24977 N24976 N24977 10
D24977 N24977 0 diode
R24978 N24977 N24978 10
D24978 N24978 0 diode
R24979 N24978 N24979 10
D24979 N24979 0 diode
R24980 N24979 N24980 10
D24980 N24980 0 diode
R24981 N24980 N24981 10
D24981 N24981 0 diode
R24982 N24981 N24982 10
D24982 N24982 0 diode
R24983 N24982 N24983 10
D24983 N24983 0 diode
R24984 N24983 N24984 10
D24984 N24984 0 diode
R24985 N24984 N24985 10
D24985 N24985 0 diode
R24986 N24985 N24986 10
D24986 N24986 0 diode
R24987 N24986 N24987 10
D24987 N24987 0 diode
R24988 N24987 N24988 10
D24988 N24988 0 diode
R24989 N24988 N24989 10
D24989 N24989 0 diode
R24990 N24989 N24990 10
D24990 N24990 0 diode
R24991 N24990 N24991 10
D24991 N24991 0 diode
R24992 N24991 N24992 10
D24992 N24992 0 diode
R24993 N24992 N24993 10
D24993 N24993 0 diode
R24994 N24993 N24994 10
D24994 N24994 0 diode
R24995 N24994 N24995 10
D24995 N24995 0 diode
R24996 N24995 N24996 10
D24996 N24996 0 diode
R24997 N24996 N24997 10
D24997 N24997 0 diode
R24998 N24997 N24998 10
D24998 N24998 0 diode
R24999 N24998 N24999 10
D24999 N24999 0 diode
R25000 N24999 N25000 10
D25000 N25000 0 diode
R25001 N25000 N25001 10
D25001 N25001 0 diode
R25002 N25001 N25002 10
D25002 N25002 0 diode
R25003 N25002 N25003 10
D25003 N25003 0 diode
R25004 N25003 N25004 10
D25004 N25004 0 diode
R25005 N25004 N25005 10
D25005 N25005 0 diode
R25006 N25005 N25006 10
D25006 N25006 0 diode
R25007 N25006 N25007 10
D25007 N25007 0 diode
R25008 N25007 N25008 10
D25008 N25008 0 diode
R25009 N25008 N25009 10
D25009 N25009 0 diode
R25010 N25009 N25010 10
D25010 N25010 0 diode
R25011 N25010 N25011 10
D25011 N25011 0 diode
R25012 N25011 N25012 10
D25012 N25012 0 diode
R25013 N25012 N25013 10
D25013 N25013 0 diode
R25014 N25013 N25014 10
D25014 N25014 0 diode
R25015 N25014 N25015 10
D25015 N25015 0 diode
R25016 N25015 N25016 10
D25016 N25016 0 diode
R25017 N25016 N25017 10
D25017 N25017 0 diode
R25018 N25017 N25018 10
D25018 N25018 0 diode
R25019 N25018 N25019 10
D25019 N25019 0 diode
R25020 N25019 N25020 10
D25020 N25020 0 diode
R25021 N25020 N25021 10
D25021 N25021 0 diode
R25022 N25021 N25022 10
D25022 N25022 0 diode
R25023 N25022 N25023 10
D25023 N25023 0 diode
R25024 N25023 N25024 10
D25024 N25024 0 diode
R25025 N25024 N25025 10
D25025 N25025 0 diode
R25026 N25025 N25026 10
D25026 N25026 0 diode
R25027 N25026 N25027 10
D25027 N25027 0 diode
R25028 N25027 N25028 10
D25028 N25028 0 diode
R25029 N25028 N25029 10
D25029 N25029 0 diode
R25030 N25029 N25030 10
D25030 N25030 0 diode
R25031 N25030 N25031 10
D25031 N25031 0 diode
R25032 N25031 N25032 10
D25032 N25032 0 diode
R25033 N25032 N25033 10
D25033 N25033 0 diode
R25034 N25033 N25034 10
D25034 N25034 0 diode
R25035 N25034 N25035 10
D25035 N25035 0 diode
R25036 N25035 N25036 10
D25036 N25036 0 diode
R25037 N25036 N25037 10
D25037 N25037 0 diode
R25038 N25037 N25038 10
D25038 N25038 0 diode
R25039 N25038 N25039 10
D25039 N25039 0 diode
R25040 N25039 N25040 10
D25040 N25040 0 diode
R25041 N25040 N25041 10
D25041 N25041 0 diode
R25042 N25041 N25042 10
D25042 N25042 0 diode
R25043 N25042 N25043 10
D25043 N25043 0 diode
R25044 N25043 N25044 10
D25044 N25044 0 diode
R25045 N25044 N25045 10
D25045 N25045 0 diode
R25046 N25045 N25046 10
D25046 N25046 0 diode
R25047 N25046 N25047 10
D25047 N25047 0 diode
R25048 N25047 N25048 10
D25048 N25048 0 diode
R25049 N25048 N25049 10
D25049 N25049 0 diode
R25050 N25049 N25050 10
D25050 N25050 0 diode
R25051 N25050 N25051 10
D25051 N25051 0 diode
R25052 N25051 N25052 10
D25052 N25052 0 diode
R25053 N25052 N25053 10
D25053 N25053 0 diode
R25054 N25053 N25054 10
D25054 N25054 0 diode
R25055 N25054 N25055 10
D25055 N25055 0 diode
R25056 N25055 N25056 10
D25056 N25056 0 diode
R25057 N25056 N25057 10
D25057 N25057 0 diode
R25058 N25057 N25058 10
D25058 N25058 0 diode
R25059 N25058 N25059 10
D25059 N25059 0 diode
R25060 N25059 N25060 10
D25060 N25060 0 diode
R25061 N25060 N25061 10
D25061 N25061 0 diode
R25062 N25061 N25062 10
D25062 N25062 0 diode
R25063 N25062 N25063 10
D25063 N25063 0 diode
R25064 N25063 N25064 10
D25064 N25064 0 diode
R25065 N25064 N25065 10
D25065 N25065 0 diode
R25066 N25065 N25066 10
D25066 N25066 0 diode
R25067 N25066 N25067 10
D25067 N25067 0 diode
R25068 N25067 N25068 10
D25068 N25068 0 diode
R25069 N25068 N25069 10
D25069 N25069 0 diode
R25070 N25069 N25070 10
D25070 N25070 0 diode
R25071 N25070 N25071 10
D25071 N25071 0 diode
R25072 N25071 N25072 10
D25072 N25072 0 diode
R25073 N25072 N25073 10
D25073 N25073 0 diode
R25074 N25073 N25074 10
D25074 N25074 0 diode
R25075 N25074 N25075 10
D25075 N25075 0 diode
R25076 N25075 N25076 10
D25076 N25076 0 diode
R25077 N25076 N25077 10
D25077 N25077 0 diode
R25078 N25077 N25078 10
D25078 N25078 0 diode
R25079 N25078 N25079 10
D25079 N25079 0 diode
R25080 N25079 N25080 10
D25080 N25080 0 diode
R25081 N25080 N25081 10
D25081 N25081 0 diode
R25082 N25081 N25082 10
D25082 N25082 0 diode
R25083 N25082 N25083 10
D25083 N25083 0 diode
R25084 N25083 N25084 10
D25084 N25084 0 diode
R25085 N25084 N25085 10
D25085 N25085 0 diode
R25086 N25085 N25086 10
D25086 N25086 0 diode
R25087 N25086 N25087 10
D25087 N25087 0 diode
R25088 N25087 N25088 10
D25088 N25088 0 diode
R25089 N25088 N25089 10
D25089 N25089 0 diode
R25090 N25089 N25090 10
D25090 N25090 0 diode
R25091 N25090 N25091 10
D25091 N25091 0 diode
R25092 N25091 N25092 10
D25092 N25092 0 diode
R25093 N25092 N25093 10
D25093 N25093 0 diode
R25094 N25093 N25094 10
D25094 N25094 0 diode
R25095 N25094 N25095 10
D25095 N25095 0 diode
R25096 N25095 N25096 10
D25096 N25096 0 diode
R25097 N25096 N25097 10
D25097 N25097 0 diode
R25098 N25097 N25098 10
D25098 N25098 0 diode
R25099 N25098 N25099 10
D25099 N25099 0 diode
R25100 N25099 N25100 10
D25100 N25100 0 diode
R25101 N25100 N25101 10
D25101 N25101 0 diode
R25102 N25101 N25102 10
D25102 N25102 0 diode
R25103 N25102 N25103 10
D25103 N25103 0 diode
R25104 N25103 N25104 10
D25104 N25104 0 diode
R25105 N25104 N25105 10
D25105 N25105 0 diode
R25106 N25105 N25106 10
D25106 N25106 0 diode
R25107 N25106 N25107 10
D25107 N25107 0 diode
R25108 N25107 N25108 10
D25108 N25108 0 diode
R25109 N25108 N25109 10
D25109 N25109 0 diode
R25110 N25109 N25110 10
D25110 N25110 0 diode
R25111 N25110 N25111 10
D25111 N25111 0 diode
R25112 N25111 N25112 10
D25112 N25112 0 diode
R25113 N25112 N25113 10
D25113 N25113 0 diode
R25114 N25113 N25114 10
D25114 N25114 0 diode
R25115 N25114 N25115 10
D25115 N25115 0 diode
R25116 N25115 N25116 10
D25116 N25116 0 diode
R25117 N25116 N25117 10
D25117 N25117 0 diode
R25118 N25117 N25118 10
D25118 N25118 0 diode
R25119 N25118 N25119 10
D25119 N25119 0 diode
R25120 N25119 N25120 10
D25120 N25120 0 diode
R25121 N25120 N25121 10
D25121 N25121 0 diode
R25122 N25121 N25122 10
D25122 N25122 0 diode
R25123 N25122 N25123 10
D25123 N25123 0 diode
R25124 N25123 N25124 10
D25124 N25124 0 diode
R25125 N25124 N25125 10
D25125 N25125 0 diode
R25126 N25125 N25126 10
D25126 N25126 0 diode
R25127 N25126 N25127 10
D25127 N25127 0 diode
R25128 N25127 N25128 10
D25128 N25128 0 diode
R25129 N25128 N25129 10
D25129 N25129 0 diode
R25130 N25129 N25130 10
D25130 N25130 0 diode
R25131 N25130 N25131 10
D25131 N25131 0 diode
R25132 N25131 N25132 10
D25132 N25132 0 diode
R25133 N25132 N25133 10
D25133 N25133 0 diode
R25134 N25133 N25134 10
D25134 N25134 0 diode
R25135 N25134 N25135 10
D25135 N25135 0 diode
R25136 N25135 N25136 10
D25136 N25136 0 diode
R25137 N25136 N25137 10
D25137 N25137 0 diode
R25138 N25137 N25138 10
D25138 N25138 0 diode
R25139 N25138 N25139 10
D25139 N25139 0 diode
R25140 N25139 N25140 10
D25140 N25140 0 diode
R25141 N25140 N25141 10
D25141 N25141 0 diode
R25142 N25141 N25142 10
D25142 N25142 0 diode
R25143 N25142 N25143 10
D25143 N25143 0 diode
R25144 N25143 N25144 10
D25144 N25144 0 diode
R25145 N25144 N25145 10
D25145 N25145 0 diode
R25146 N25145 N25146 10
D25146 N25146 0 diode
R25147 N25146 N25147 10
D25147 N25147 0 diode
R25148 N25147 N25148 10
D25148 N25148 0 diode
R25149 N25148 N25149 10
D25149 N25149 0 diode
R25150 N25149 N25150 10
D25150 N25150 0 diode
R25151 N25150 N25151 10
D25151 N25151 0 diode
R25152 N25151 N25152 10
D25152 N25152 0 diode
R25153 N25152 N25153 10
D25153 N25153 0 diode
R25154 N25153 N25154 10
D25154 N25154 0 diode
R25155 N25154 N25155 10
D25155 N25155 0 diode
R25156 N25155 N25156 10
D25156 N25156 0 diode
R25157 N25156 N25157 10
D25157 N25157 0 diode
R25158 N25157 N25158 10
D25158 N25158 0 diode
R25159 N25158 N25159 10
D25159 N25159 0 diode
R25160 N25159 N25160 10
D25160 N25160 0 diode
R25161 N25160 N25161 10
D25161 N25161 0 diode
R25162 N25161 N25162 10
D25162 N25162 0 diode
R25163 N25162 N25163 10
D25163 N25163 0 diode
R25164 N25163 N25164 10
D25164 N25164 0 diode
R25165 N25164 N25165 10
D25165 N25165 0 diode
R25166 N25165 N25166 10
D25166 N25166 0 diode
R25167 N25166 N25167 10
D25167 N25167 0 diode
R25168 N25167 N25168 10
D25168 N25168 0 diode
R25169 N25168 N25169 10
D25169 N25169 0 diode
R25170 N25169 N25170 10
D25170 N25170 0 diode
R25171 N25170 N25171 10
D25171 N25171 0 diode
R25172 N25171 N25172 10
D25172 N25172 0 diode
R25173 N25172 N25173 10
D25173 N25173 0 diode
R25174 N25173 N25174 10
D25174 N25174 0 diode
R25175 N25174 N25175 10
D25175 N25175 0 diode
R25176 N25175 N25176 10
D25176 N25176 0 diode
R25177 N25176 N25177 10
D25177 N25177 0 diode
R25178 N25177 N25178 10
D25178 N25178 0 diode
R25179 N25178 N25179 10
D25179 N25179 0 diode
R25180 N25179 N25180 10
D25180 N25180 0 diode
R25181 N25180 N25181 10
D25181 N25181 0 diode
R25182 N25181 N25182 10
D25182 N25182 0 diode
R25183 N25182 N25183 10
D25183 N25183 0 diode
R25184 N25183 N25184 10
D25184 N25184 0 diode
R25185 N25184 N25185 10
D25185 N25185 0 diode
R25186 N25185 N25186 10
D25186 N25186 0 diode
R25187 N25186 N25187 10
D25187 N25187 0 diode
R25188 N25187 N25188 10
D25188 N25188 0 diode
R25189 N25188 N25189 10
D25189 N25189 0 diode
R25190 N25189 N25190 10
D25190 N25190 0 diode
R25191 N25190 N25191 10
D25191 N25191 0 diode
R25192 N25191 N25192 10
D25192 N25192 0 diode
R25193 N25192 N25193 10
D25193 N25193 0 diode
R25194 N25193 N25194 10
D25194 N25194 0 diode
R25195 N25194 N25195 10
D25195 N25195 0 diode
R25196 N25195 N25196 10
D25196 N25196 0 diode
R25197 N25196 N25197 10
D25197 N25197 0 diode
R25198 N25197 N25198 10
D25198 N25198 0 diode
R25199 N25198 N25199 10
D25199 N25199 0 diode
R25200 N25199 N25200 10
D25200 N25200 0 diode
R25201 N25200 N25201 10
D25201 N25201 0 diode
R25202 N25201 N25202 10
D25202 N25202 0 diode
R25203 N25202 N25203 10
D25203 N25203 0 diode
R25204 N25203 N25204 10
D25204 N25204 0 diode
R25205 N25204 N25205 10
D25205 N25205 0 diode
R25206 N25205 N25206 10
D25206 N25206 0 diode
R25207 N25206 N25207 10
D25207 N25207 0 diode
R25208 N25207 N25208 10
D25208 N25208 0 diode
R25209 N25208 N25209 10
D25209 N25209 0 diode
R25210 N25209 N25210 10
D25210 N25210 0 diode
R25211 N25210 N25211 10
D25211 N25211 0 diode
R25212 N25211 N25212 10
D25212 N25212 0 diode
R25213 N25212 N25213 10
D25213 N25213 0 diode
R25214 N25213 N25214 10
D25214 N25214 0 diode
R25215 N25214 N25215 10
D25215 N25215 0 diode
R25216 N25215 N25216 10
D25216 N25216 0 diode
R25217 N25216 N25217 10
D25217 N25217 0 diode
R25218 N25217 N25218 10
D25218 N25218 0 diode
R25219 N25218 N25219 10
D25219 N25219 0 diode
R25220 N25219 N25220 10
D25220 N25220 0 diode
R25221 N25220 N25221 10
D25221 N25221 0 diode
R25222 N25221 N25222 10
D25222 N25222 0 diode
R25223 N25222 N25223 10
D25223 N25223 0 diode
R25224 N25223 N25224 10
D25224 N25224 0 diode
R25225 N25224 N25225 10
D25225 N25225 0 diode
R25226 N25225 N25226 10
D25226 N25226 0 diode
R25227 N25226 N25227 10
D25227 N25227 0 diode
R25228 N25227 N25228 10
D25228 N25228 0 diode
R25229 N25228 N25229 10
D25229 N25229 0 diode
R25230 N25229 N25230 10
D25230 N25230 0 diode
R25231 N25230 N25231 10
D25231 N25231 0 diode
R25232 N25231 N25232 10
D25232 N25232 0 diode
R25233 N25232 N25233 10
D25233 N25233 0 diode
R25234 N25233 N25234 10
D25234 N25234 0 diode
R25235 N25234 N25235 10
D25235 N25235 0 diode
R25236 N25235 N25236 10
D25236 N25236 0 diode
R25237 N25236 N25237 10
D25237 N25237 0 diode
R25238 N25237 N25238 10
D25238 N25238 0 diode
R25239 N25238 N25239 10
D25239 N25239 0 diode
R25240 N25239 N25240 10
D25240 N25240 0 diode
R25241 N25240 N25241 10
D25241 N25241 0 diode
R25242 N25241 N25242 10
D25242 N25242 0 diode
R25243 N25242 N25243 10
D25243 N25243 0 diode
R25244 N25243 N25244 10
D25244 N25244 0 diode
R25245 N25244 N25245 10
D25245 N25245 0 diode
R25246 N25245 N25246 10
D25246 N25246 0 diode
R25247 N25246 N25247 10
D25247 N25247 0 diode
R25248 N25247 N25248 10
D25248 N25248 0 diode
R25249 N25248 N25249 10
D25249 N25249 0 diode
R25250 N25249 N25250 10
D25250 N25250 0 diode
R25251 N25250 N25251 10
D25251 N25251 0 diode
R25252 N25251 N25252 10
D25252 N25252 0 diode
R25253 N25252 N25253 10
D25253 N25253 0 diode
R25254 N25253 N25254 10
D25254 N25254 0 diode
R25255 N25254 N25255 10
D25255 N25255 0 diode
R25256 N25255 N25256 10
D25256 N25256 0 diode
R25257 N25256 N25257 10
D25257 N25257 0 diode
R25258 N25257 N25258 10
D25258 N25258 0 diode
R25259 N25258 N25259 10
D25259 N25259 0 diode
R25260 N25259 N25260 10
D25260 N25260 0 diode
R25261 N25260 N25261 10
D25261 N25261 0 diode
R25262 N25261 N25262 10
D25262 N25262 0 diode
R25263 N25262 N25263 10
D25263 N25263 0 diode
R25264 N25263 N25264 10
D25264 N25264 0 diode
R25265 N25264 N25265 10
D25265 N25265 0 diode
R25266 N25265 N25266 10
D25266 N25266 0 diode
R25267 N25266 N25267 10
D25267 N25267 0 diode
R25268 N25267 N25268 10
D25268 N25268 0 diode
R25269 N25268 N25269 10
D25269 N25269 0 diode
R25270 N25269 N25270 10
D25270 N25270 0 diode
R25271 N25270 N25271 10
D25271 N25271 0 diode
R25272 N25271 N25272 10
D25272 N25272 0 diode
R25273 N25272 N25273 10
D25273 N25273 0 diode
R25274 N25273 N25274 10
D25274 N25274 0 diode
R25275 N25274 N25275 10
D25275 N25275 0 diode
R25276 N25275 N25276 10
D25276 N25276 0 diode
R25277 N25276 N25277 10
D25277 N25277 0 diode
R25278 N25277 N25278 10
D25278 N25278 0 diode
R25279 N25278 N25279 10
D25279 N25279 0 diode
R25280 N25279 N25280 10
D25280 N25280 0 diode
R25281 N25280 N25281 10
D25281 N25281 0 diode
R25282 N25281 N25282 10
D25282 N25282 0 diode
R25283 N25282 N25283 10
D25283 N25283 0 diode
R25284 N25283 N25284 10
D25284 N25284 0 diode
R25285 N25284 N25285 10
D25285 N25285 0 diode
R25286 N25285 N25286 10
D25286 N25286 0 diode
R25287 N25286 N25287 10
D25287 N25287 0 diode
R25288 N25287 N25288 10
D25288 N25288 0 diode
R25289 N25288 N25289 10
D25289 N25289 0 diode
R25290 N25289 N25290 10
D25290 N25290 0 diode
R25291 N25290 N25291 10
D25291 N25291 0 diode
R25292 N25291 N25292 10
D25292 N25292 0 diode
R25293 N25292 N25293 10
D25293 N25293 0 diode
R25294 N25293 N25294 10
D25294 N25294 0 diode
R25295 N25294 N25295 10
D25295 N25295 0 diode
R25296 N25295 N25296 10
D25296 N25296 0 diode
R25297 N25296 N25297 10
D25297 N25297 0 diode
R25298 N25297 N25298 10
D25298 N25298 0 diode
R25299 N25298 N25299 10
D25299 N25299 0 diode
R25300 N25299 N25300 10
D25300 N25300 0 diode
R25301 N25300 N25301 10
D25301 N25301 0 diode
R25302 N25301 N25302 10
D25302 N25302 0 diode
R25303 N25302 N25303 10
D25303 N25303 0 diode
R25304 N25303 N25304 10
D25304 N25304 0 diode
R25305 N25304 N25305 10
D25305 N25305 0 diode
R25306 N25305 N25306 10
D25306 N25306 0 diode
R25307 N25306 N25307 10
D25307 N25307 0 diode
R25308 N25307 N25308 10
D25308 N25308 0 diode
R25309 N25308 N25309 10
D25309 N25309 0 diode
R25310 N25309 N25310 10
D25310 N25310 0 diode
R25311 N25310 N25311 10
D25311 N25311 0 diode
R25312 N25311 N25312 10
D25312 N25312 0 diode
R25313 N25312 N25313 10
D25313 N25313 0 diode
R25314 N25313 N25314 10
D25314 N25314 0 diode
R25315 N25314 N25315 10
D25315 N25315 0 diode
R25316 N25315 N25316 10
D25316 N25316 0 diode
R25317 N25316 N25317 10
D25317 N25317 0 diode
R25318 N25317 N25318 10
D25318 N25318 0 diode
R25319 N25318 N25319 10
D25319 N25319 0 diode
R25320 N25319 N25320 10
D25320 N25320 0 diode
R25321 N25320 N25321 10
D25321 N25321 0 diode
R25322 N25321 N25322 10
D25322 N25322 0 diode
R25323 N25322 N25323 10
D25323 N25323 0 diode
R25324 N25323 N25324 10
D25324 N25324 0 diode
R25325 N25324 N25325 10
D25325 N25325 0 diode
R25326 N25325 N25326 10
D25326 N25326 0 diode
R25327 N25326 N25327 10
D25327 N25327 0 diode
R25328 N25327 N25328 10
D25328 N25328 0 diode
R25329 N25328 N25329 10
D25329 N25329 0 diode
R25330 N25329 N25330 10
D25330 N25330 0 diode
R25331 N25330 N25331 10
D25331 N25331 0 diode
R25332 N25331 N25332 10
D25332 N25332 0 diode
R25333 N25332 N25333 10
D25333 N25333 0 diode
R25334 N25333 N25334 10
D25334 N25334 0 diode
R25335 N25334 N25335 10
D25335 N25335 0 diode
R25336 N25335 N25336 10
D25336 N25336 0 diode
R25337 N25336 N25337 10
D25337 N25337 0 diode
R25338 N25337 N25338 10
D25338 N25338 0 diode
R25339 N25338 N25339 10
D25339 N25339 0 diode
R25340 N25339 N25340 10
D25340 N25340 0 diode
R25341 N25340 N25341 10
D25341 N25341 0 diode
R25342 N25341 N25342 10
D25342 N25342 0 diode
R25343 N25342 N25343 10
D25343 N25343 0 diode
R25344 N25343 N25344 10
D25344 N25344 0 diode
R25345 N25344 N25345 10
D25345 N25345 0 diode
R25346 N25345 N25346 10
D25346 N25346 0 diode
R25347 N25346 N25347 10
D25347 N25347 0 diode
R25348 N25347 N25348 10
D25348 N25348 0 diode
R25349 N25348 N25349 10
D25349 N25349 0 diode
R25350 N25349 N25350 10
D25350 N25350 0 diode
R25351 N25350 N25351 10
D25351 N25351 0 diode
R25352 N25351 N25352 10
D25352 N25352 0 diode
R25353 N25352 N25353 10
D25353 N25353 0 diode
R25354 N25353 N25354 10
D25354 N25354 0 diode
R25355 N25354 N25355 10
D25355 N25355 0 diode
R25356 N25355 N25356 10
D25356 N25356 0 diode
R25357 N25356 N25357 10
D25357 N25357 0 diode
R25358 N25357 N25358 10
D25358 N25358 0 diode
R25359 N25358 N25359 10
D25359 N25359 0 diode
R25360 N25359 N25360 10
D25360 N25360 0 diode
R25361 N25360 N25361 10
D25361 N25361 0 diode
R25362 N25361 N25362 10
D25362 N25362 0 diode
R25363 N25362 N25363 10
D25363 N25363 0 diode
R25364 N25363 N25364 10
D25364 N25364 0 diode
R25365 N25364 N25365 10
D25365 N25365 0 diode
R25366 N25365 N25366 10
D25366 N25366 0 diode
R25367 N25366 N25367 10
D25367 N25367 0 diode
R25368 N25367 N25368 10
D25368 N25368 0 diode
R25369 N25368 N25369 10
D25369 N25369 0 diode
R25370 N25369 N25370 10
D25370 N25370 0 diode
R25371 N25370 N25371 10
D25371 N25371 0 diode
R25372 N25371 N25372 10
D25372 N25372 0 diode
R25373 N25372 N25373 10
D25373 N25373 0 diode
R25374 N25373 N25374 10
D25374 N25374 0 diode
R25375 N25374 N25375 10
D25375 N25375 0 diode
R25376 N25375 N25376 10
D25376 N25376 0 diode
R25377 N25376 N25377 10
D25377 N25377 0 diode
R25378 N25377 N25378 10
D25378 N25378 0 diode
R25379 N25378 N25379 10
D25379 N25379 0 diode
R25380 N25379 N25380 10
D25380 N25380 0 diode
R25381 N25380 N25381 10
D25381 N25381 0 diode
R25382 N25381 N25382 10
D25382 N25382 0 diode
R25383 N25382 N25383 10
D25383 N25383 0 diode
R25384 N25383 N25384 10
D25384 N25384 0 diode
R25385 N25384 N25385 10
D25385 N25385 0 diode
R25386 N25385 N25386 10
D25386 N25386 0 diode
R25387 N25386 N25387 10
D25387 N25387 0 diode
R25388 N25387 N25388 10
D25388 N25388 0 diode
R25389 N25388 N25389 10
D25389 N25389 0 diode
R25390 N25389 N25390 10
D25390 N25390 0 diode
R25391 N25390 N25391 10
D25391 N25391 0 diode
R25392 N25391 N25392 10
D25392 N25392 0 diode
R25393 N25392 N25393 10
D25393 N25393 0 diode
R25394 N25393 N25394 10
D25394 N25394 0 diode
R25395 N25394 N25395 10
D25395 N25395 0 diode
R25396 N25395 N25396 10
D25396 N25396 0 diode
R25397 N25396 N25397 10
D25397 N25397 0 diode
R25398 N25397 N25398 10
D25398 N25398 0 diode
R25399 N25398 N25399 10
D25399 N25399 0 diode
R25400 N25399 N25400 10
D25400 N25400 0 diode
R25401 N25400 N25401 10
D25401 N25401 0 diode
R25402 N25401 N25402 10
D25402 N25402 0 diode
R25403 N25402 N25403 10
D25403 N25403 0 diode
R25404 N25403 N25404 10
D25404 N25404 0 diode
R25405 N25404 N25405 10
D25405 N25405 0 diode
R25406 N25405 N25406 10
D25406 N25406 0 diode
R25407 N25406 N25407 10
D25407 N25407 0 diode
R25408 N25407 N25408 10
D25408 N25408 0 diode
R25409 N25408 N25409 10
D25409 N25409 0 diode
R25410 N25409 N25410 10
D25410 N25410 0 diode
R25411 N25410 N25411 10
D25411 N25411 0 diode
R25412 N25411 N25412 10
D25412 N25412 0 diode
R25413 N25412 N25413 10
D25413 N25413 0 diode
R25414 N25413 N25414 10
D25414 N25414 0 diode
R25415 N25414 N25415 10
D25415 N25415 0 diode
R25416 N25415 N25416 10
D25416 N25416 0 diode
R25417 N25416 N25417 10
D25417 N25417 0 diode
R25418 N25417 N25418 10
D25418 N25418 0 diode
R25419 N25418 N25419 10
D25419 N25419 0 diode
R25420 N25419 N25420 10
D25420 N25420 0 diode
R25421 N25420 N25421 10
D25421 N25421 0 diode
R25422 N25421 N25422 10
D25422 N25422 0 diode
R25423 N25422 N25423 10
D25423 N25423 0 diode
R25424 N25423 N25424 10
D25424 N25424 0 diode
R25425 N25424 N25425 10
D25425 N25425 0 diode
R25426 N25425 N25426 10
D25426 N25426 0 diode
R25427 N25426 N25427 10
D25427 N25427 0 diode
R25428 N25427 N25428 10
D25428 N25428 0 diode
R25429 N25428 N25429 10
D25429 N25429 0 diode
R25430 N25429 N25430 10
D25430 N25430 0 diode
R25431 N25430 N25431 10
D25431 N25431 0 diode
R25432 N25431 N25432 10
D25432 N25432 0 diode
R25433 N25432 N25433 10
D25433 N25433 0 diode
R25434 N25433 N25434 10
D25434 N25434 0 diode
R25435 N25434 N25435 10
D25435 N25435 0 diode
R25436 N25435 N25436 10
D25436 N25436 0 diode
R25437 N25436 N25437 10
D25437 N25437 0 diode
R25438 N25437 N25438 10
D25438 N25438 0 diode
R25439 N25438 N25439 10
D25439 N25439 0 diode
R25440 N25439 N25440 10
D25440 N25440 0 diode
R25441 N25440 N25441 10
D25441 N25441 0 diode
R25442 N25441 N25442 10
D25442 N25442 0 diode
R25443 N25442 N25443 10
D25443 N25443 0 diode
R25444 N25443 N25444 10
D25444 N25444 0 diode
R25445 N25444 N25445 10
D25445 N25445 0 diode
R25446 N25445 N25446 10
D25446 N25446 0 diode
R25447 N25446 N25447 10
D25447 N25447 0 diode
R25448 N25447 N25448 10
D25448 N25448 0 diode
R25449 N25448 N25449 10
D25449 N25449 0 diode
R25450 N25449 N25450 10
D25450 N25450 0 diode
R25451 N25450 N25451 10
D25451 N25451 0 diode
R25452 N25451 N25452 10
D25452 N25452 0 diode
R25453 N25452 N25453 10
D25453 N25453 0 diode
R25454 N25453 N25454 10
D25454 N25454 0 diode
R25455 N25454 N25455 10
D25455 N25455 0 diode
R25456 N25455 N25456 10
D25456 N25456 0 diode
R25457 N25456 N25457 10
D25457 N25457 0 diode
R25458 N25457 N25458 10
D25458 N25458 0 diode
R25459 N25458 N25459 10
D25459 N25459 0 diode
R25460 N25459 N25460 10
D25460 N25460 0 diode
R25461 N25460 N25461 10
D25461 N25461 0 diode
R25462 N25461 N25462 10
D25462 N25462 0 diode
R25463 N25462 N25463 10
D25463 N25463 0 diode
R25464 N25463 N25464 10
D25464 N25464 0 diode
R25465 N25464 N25465 10
D25465 N25465 0 diode
R25466 N25465 N25466 10
D25466 N25466 0 diode
R25467 N25466 N25467 10
D25467 N25467 0 diode
R25468 N25467 N25468 10
D25468 N25468 0 diode
R25469 N25468 N25469 10
D25469 N25469 0 diode
R25470 N25469 N25470 10
D25470 N25470 0 diode
R25471 N25470 N25471 10
D25471 N25471 0 diode
R25472 N25471 N25472 10
D25472 N25472 0 diode
R25473 N25472 N25473 10
D25473 N25473 0 diode
R25474 N25473 N25474 10
D25474 N25474 0 diode
R25475 N25474 N25475 10
D25475 N25475 0 diode
R25476 N25475 N25476 10
D25476 N25476 0 diode
R25477 N25476 N25477 10
D25477 N25477 0 diode
R25478 N25477 N25478 10
D25478 N25478 0 diode
R25479 N25478 N25479 10
D25479 N25479 0 diode
R25480 N25479 N25480 10
D25480 N25480 0 diode
R25481 N25480 N25481 10
D25481 N25481 0 diode
R25482 N25481 N25482 10
D25482 N25482 0 diode
R25483 N25482 N25483 10
D25483 N25483 0 diode
R25484 N25483 N25484 10
D25484 N25484 0 diode
R25485 N25484 N25485 10
D25485 N25485 0 diode
R25486 N25485 N25486 10
D25486 N25486 0 diode
R25487 N25486 N25487 10
D25487 N25487 0 diode
R25488 N25487 N25488 10
D25488 N25488 0 diode
R25489 N25488 N25489 10
D25489 N25489 0 diode
R25490 N25489 N25490 10
D25490 N25490 0 diode
R25491 N25490 N25491 10
D25491 N25491 0 diode
R25492 N25491 N25492 10
D25492 N25492 0 diode
R25493 N25492 N25493 10
D25493 N25493 0 diode
R25494 N25493 N25494 10
D25494 N25494 0 diode
R25495 N25494 N25495 10
D25495 N25495 0 diode
R25496 N25495 N25496 10
D25496 N25496 0 diode
R25497 N25496 N25497 10
D25497 N25497 0 diode
R25498 N25497 N25498 10
D25498 N25498 0 diode
R25499 N25498 N25499 10
D25499 N25499 0 diode
R25500 N25499 N25500 10
D25500 N25500 0 diode
R25501 N25500 N25501 10
D25501 N25501 0 diode
R25502 N25501 N25502 10
D25502 N25502 0 diode
R25503 N25502 N25503 10
D25503 N25503 0 diode
R25504 N25503 N25504 10
D25504 N25504 0 diode
R25505 N25504 N25505 10
D25505 N25505 0 diode
R25506 N25505 N25506 10
D25506 N25506 0 diode
R25507 N25506 N25507 10
D25507 N25507 0 diode
R25508 N25507 N25508 10
D25508 N25508 0 diode
R25509 N25508 N25509 10
D25509 N25509 0 diode
R25510 N25509 N25510 10
D25510 N25510 0 diode
R25511 N25510 N25511 10
D25511 N25511 0 diode
R25512 N25511 N25512 10
D25512 N25512 0 diode
R25513 N25512 N25513 10
D25513 N25513 0 diode
R25514 N25513 N25514 10
D25514 N25514 0 diode
R25515 N25514 N25515 10
D25515 N25515 0 diode
R25516 N25515 N25516 10
D25516 N25516 0 diode
R25517 N25516 N25517 10
D25517 N25517 0 diode
R25518 N25517 N25518 10
D25518 N25518 0 diode
R25519 N25518 N25519 10
D25519 N25519 0 diode
R25520 N25519 N25520 10
D25520 N25520 0 diode
R25521 N25520 N25521 10
D25521 N25521 0 diode
R25522 N25521 N25522 10
D25522 N25522 0 diode
R25523 N25522 N25523 10
D25523 N25523 0 diode
R25524 N25523 N25524 10
D25524 N25524 0 diode
R25525 N25524 N25525 10
D25525 N25525 0 diode
R25526 N25525 N25526 10
D25526 N25526 0 diode
R25527 N25526 N25527 10
D25527 N25527 0 diode
R25528 N25527 N25528 10
D25528 N25528 0 diode
R25529 N25528 N25529 10
D25529 N25529 0 diode
R25530 N25529 N25530 10
D25530 N25530 0 diode
R25531 N25530 N25531 10
D25531 N25531 0 diode
R25532 N25531 N25532 10
D25532 N25532 0 diode
R25533 N25532 N25533 10
D25533 N25533 0 diode
R25534 N25533 N25534 10
D25534 N25534 0 diode
R25535 N25534 N25535 10
D25535 N25535 0 diode
R25536 N25535 N25536 10
D25536 N25536 0 diode
R25537 N25536 N25537 10
D25537 N25537 0 diode
R25538 N25537 N25538 10
D25538 N25538 0 diode
R25539 N25538 N25539 10
D25539 N25539 0 diode
R25540 N25539 N25540 10
D25540 N25540 0 diode
R25541 N25540 N25541 10
D25541 N25541 0 diode
R25542 N25541 N25542 10
D25542 N25542 0 diode
R25543 N25542 N25543 10
D25543 N25543 0 diode
R25544 N25543 N25544 10
D25544 N25544 0 diode
R25545 N25544 N25545 10
D25545 N25545 0 diode
R25546 N25545 N25546 10
D25546 N25546 0 diode
R25547 N25546 N25547 10
D25547 N25547 0 diode
R25548 N25547 N25548 10
D25548 N25548 0 diode
R25549 N25548 N25549 10
D25549 N25549 0 diode
R25550 N25549 N25550 10
D25550 N25550 0 diode
R25551 N25550 N25551 10
D25551 N25551 0 diode
R25552 N25551 N25552 10
D25552 N25552 0 diode
R25553 N25552 N25553 10
D25553 N25553 0 diode
R25554 N25553 N25554 10
D25554 N25554 0 diode
R25555 N25554 N25555 10
D25555 N25555 0 diode
R25556 N25555 N25556 10
D25556 N25556 0 diode
R25557 N25556 N25557 10
D25557 N25557 0 diode
R25558 N25557 N25558 10
D25558 N25558 0 diode
R25559 N25558 N25559 10
D25559 N25559 0 diode
R25560 N25559 N25560 10
D25560 N25560 0 diode
R25561 N25560 N25561 10
D25561 N25561 0 diode
R25562 N25561 N25562 10
D25562 N25562 0 diode
R25563 N25562 N25563 10
D25563 N25563 0 diode
R25564 N25563 N25564 10
D25564 N25564 0 diode
R25565 N25564 N25565 10
D25565 N25565 0 diode
R25566 N25565 N25566 10
D25566 N25566 0 diode
R25567 N25566 N25567 10
D25567 N25567 0 diode
R25568 N25567 N25568 10
D25568 N25568 0 diode
R25569 N25568 N25569 10
D25569 N25569 0 diode
R25570 N25569 N25570 10
D25570 N25570 0 diode
R25571 N25570 N25571 10
D25571 N25571 0 diode
R25572 N25571 N25572 10
D25572 N25572 0 diode
R25573 N25572 N25573 10
D25573 N25573 0 diode
R25574 N25573 N25574 10
D25574 N25574 0 diode
R25575 N25574 N25575 10
D25575 N25575 0 diode
R25576 N25575 N25576 10
D25576 N25576 0 diode
R25577 N25576 N25577 10
D25577 N25577 0 diode
R25578 N25577 N25578 10
D25578 N25578 0 diode
R25579 N25578 N25579 10
D25579 N25579 0 diode
R25580 N25579 N25580 10
D25580 N25580 0 diode
R25581 N25580 N25581 10
D25581 N25581 0 diode
R25582 N25581 N25582 10
D25582 N25582 0 diode
R25583 N25582 N25583 10
D25583 N25583 0 diode
R25584 N25583 N25584 10
D25584 N25584 0 diode
R25585 N25584 N25585 10
D25585 N25585 0 diode
R25586 N25585 N25586 10
D25586 N25586 0 diode
R25587 N25586 N25587 10
D25587 N25587 0 diode
R25588 N25587 N25588 10
D25588 N25588 0 diode
R25589 N25588 N25589 10
D25589 N25589 0 diode
R25590 N25589 N25590 10
D25590 N25590 0 diode
R25591 N25590 N25591 10
D25591 N25591 0 diode
R25592 N25591 N25592 10
D25592 N25592 0 diode
R25593 N25592 N25593 10
D25593 N25593 0 diode
R25594 N25593 N25594 10
D25594 N25594 0 diode
R25595 N25594 N25595 10
D25595 N25595 0 diode
R25596 N25595 N25596 10
D25596 N25596 0 diode
R25597 N25596 N25597 10
D25597 N25597 0 diode
R25598 N25597 N25598 10
D25598 N25598 0 diode
R25599 N25598 N25599 10
D25599 N25599 0 diode
R25600 N25599 N25600 10
D25600 N25600 0 diode
R25601 N25600 N25601 10
D25601 N25601 0 diode
R25602 N25601 N25602 10
D25602 N25602 0 diode
R25603 N25602 N25603 10
D25603 N25603 0 diode
R25604 N25603 N25604 10
D25604 N25604 0 diode
R25605 N25604 N25605 10
D25605 N25605 0 diode
R25606 N25605 N25606 10
D25606 N25606 0 diode
R25607 N25606 N25607 10
D25607 N25607 0 diode
R25608 N25607 N25608 10
D25608 N25608 0 diode
R25609 N25608 N25609 10
D25609 N25609 0 diode
R25610 N25609 N25610 10
D25610 N25610 0 diode
R25611 N25610 N25611 10
D25611 N25611 0 diode
R25612 N25611 N25612 10
D25612 N25612 0 diode
R25613 N25612 N25613 10
D25613 N25613 0 diode
R25614 N25613 N25614 10
D25614 N25614 0 diode
R25615 N25614 N25615 10
D25615 N25615 0 diode
R25616 N25615 N25616 10
D25616 N25616 0 diode
R25617 N25616 N25617 10
D25617 N25617 0 diode
R25618 N25617 N25618 10
D25618 N25618 0 diode
R25619 N25618 N25619 10
D25619 N25619 0 diode
R25620 N25619 N25620 10
D25620 N25620 0 diode
R25621 N25620 N25621 10
D25621 N25621 0 diode
R25622 N25621 N25622 10
D25622 N25622 0 diode
R25623 N25622 N25623 10
D25623 N25623 0 diode
R25624 N25623 N25624 10
D25624 N25624 0 diode
R25625 N25624 N25625 10
D25625 N25625 0 diode
R25626 N25625 N25626 10
D25626 N25626 0 diode
R25627 N25626 N25627 10
D25627 N25627 0 diode
R25628 N25627 N25628 10
D25628 N25628 0 diode
R25629 N25628 N25629 10
D25629 N25629 0 diode
R25630 N25629 N25630 10
D25630 N25630 0 diode
R25631 N25630 N25631 10
D25631 N25631 0 diode
R25632 N25631 N25632 10
D25632 N25632 0 diode
R25633 N25632 N25633 10
D25633 N25633 0 diode
R25634 N25633 N25634 10
D25634 N25634 0 diode
R25635 N25634 N25635 10
D25635 N25635 0 diode
R25636 N25635 N25636 10
D25636 N25636 0 diode
R25637 N25636 N25637 10
D25637 N25637 0 diode
R25638 N25637 N25638 10
D25638 N25638 0 diode
R25639 N25638 N25639 10
D25639 N25639 0 diode
R25640 N25639 N25640 10
D25640 N25640 0 diode
R25641 N25640 N25641 10
D25641 N25641 0 diode
R25642 N25641 N25642 10
D25642 N25642 0 diode
R25643 N25642 N25643 10
D25643 N25643 0 diode
R25644 N25643 N25644 10
D25644 N25644 0 diode
R25645 N25644 N25645 10
D25645 N25645 0 diode
R25646 N25645 N25646 10
D25646 N25646 0 diode
R25647 N25646 N25647 10
D25647 N25647 0 diode
R25648 N25647 N25648 10
D25648 N25648 0 diode
R25649 N25648 N25649 10
D25649 N25649 0 diode
R25650 N25649 N25650 10
D25650 N25650 0 diode
R25651 N25650 N25651 10
D25651 N25651 0 diode
R25652 N25651 N25652 10
D25652 N25652 0 diode
R25653 N25652 N25653 10
D25653 N25653 0 diode
R25654 N25653 N25654 10
D25654 N25654 0 diode
R25655 N25654 N25655 10
D25655 N25655 0 diode
R25656 N25655 N25656 10
D25656 N25656 0 diode
R25657 N25656 N25657 10
D25657 N25657 0 diode
R25658 N25657 N25658 10
D25658 N25658 0 diode
R25659 N25658 N25659 10
D25659 N25659 0 diode
R25660 N25659 N25660 10
D25660 N25660 0 diode
R25661 N25660 N25661 10
D25661 N25661 0 diode
R25662 N25661 N25662 10
D25662 N25662 0 diode
R25663 N25662 N25663 10
D25663 N25663 0 diode
R25664 N25663 N25664 10
D25664 N25664 0 diode
R25665 N25664 N25665 10
D25665 N25665 0 diode
R25666 N25665 N25666 10
D25666 N25666 0 diode
R25667 N25666 N25667 10
D25667 N25667 0 diode
R25668 N25667 N25668 10
D25668 N25668 0 diode
R25669 N25668 N25669 10
D25669 N25669 0 diode
R25670 N25669 N25670 10
D25670 N25670 0 diode
R25671 N25670 N25671 10
D25671 N25671 0 diode
R25672 N25671 N25672 10
D25672 N25672 0 diode
R25673 N25672 N25673 10
D25673 N25673 0 diode
R25674 N25673 N25674 10
D25674 N25674 0 diode
R25675 N25674 N25675 10
D25675 N25675 0 diode
R25676 N25675 N25676 10
D25676 N25676 0 diode
R25677 N25676 N25677 10
D25677 N25677 0 diode
R25678 N25677 N25678 10
D25678 N25678 0 diode
R25679 N25678 N25679 10
D25679 N25679 0 diode
R25680 N25679 N25680 10
D25680 N25680 0 diode
R25681 N25680 N25681 10
D25681 N25681 0 diode
R25682 N25681 N25682 10
D25682 N25682 0 diode
R25683 N25682 N25683 10
D25683 N25683 0 diode
R25684 N25683 N25684 10
D25684 N25684 0 diode
R25685 N25684 N25685 10
D25685 N25685 0 diode
R25686 N25685 N25686 10
D25686 N25686 0 diode
R25687 N25686 N25687 10
D25687 N25687 0 diode
R25688 N25687 N25688 10
D25688 N25688 0 diode
R25689 N25688 N25689 10
D25689 N25689 0 diode
R25690 N25689 N25690 10
D25690 N25690 0 diode
R25691 N25690 N25691 10
D25691 N25691 0 diode
R25692 N25691 N25692 10
D25692 N25692 0 diode
R25693 N25692 N25693 10
D25693 N25693 0 diode
R25694 N25693 N25694 10
D25694 N25694 0 diode
R25695 N25694 N25695 10
D25695 N25695 0 diode
R25696 N25695 N25696 10
D25696 N25696 0 diode
R25697 N25696 N25697 10
D25697 N25697 0 diode
R25698 N25697 N25698 10
D25698 N25698 0 diode
R25699 N25698 N25699 10
D25699 N25699 0 diode
R25700 N25699 N25700 10
D25700 N25700 0 diode
R25701 N25700 N25701 10
D25701 N25701 0 diode
R25702 N25701 N25702 10
D25702 N25702 0 diode
R25703 N25702 N25703 10
D25703 N25703 0 diode
R25704 N25703 N25704 10
D25704 N25704 0 diode
R25705 N25704 N25705 10
D25705 N25705 0 diode
R25706 N25705 N25706 10
D25706 N25706 0 diode
R25707 N25706 N25707 10
D25707 N25707 0 diode
R25708 N25707 N25708 10
D25708 N25708 0 diode
R25709 N25708 N25709 10
D25709 N25709 0 diode
R25710 N25709 N25710 10
D25710 N25710 0 diode
R25711 N25710 N25711 10
D25711 N25711 0 diode
R25712 N25711 N25712 10
D25712 N25712 0 diode
R25713 N25712 N25713 10
D25713 N25713 0 diode
R25714 N25713 N25714 10
D25714 N25714 0 diode
R25715 N25714 N25715 10
D25715 N25715 0 diode
R25716 N25715 N25716 10
D25716 N25716 0 diode
R25717 N25716 N25717 10
D25717 N25717 0 diode
R25718 N25717 N25718 10
D25718 N25718 0 diode
R25719 N25718 N25719 10
D25719 N25719 0 diode
R25720 N25719 N25720 10
D25720 N25720 0 diode
R25721 N25720 N25721 10
D25721 N25721 0 diode
R25722 N25721 N25722 10
D25722 N25722 0 diode
R25723 N25722 N25723 10
D25723 N25723 0 diode
R25724 N25723 N25724 10
D25724 N25724 0 diode
R25725 N25724 N25725 10
D25725 N25725 0 diode
R25726 N25725 N25726 10
D25726 N25726 0 diode
R25727 N25726 N25727 10
D25727 N25727 0 diode
R25728 N25727 N25728 10
D25728 N25728 0 diode
R25729 N25728 N25729 10
D25729 N25729 0 diode
R25730 N25729 N25730 10
D25730 N25730 0 diode
R25731 N25730 N25731 10
D25731 N25731 0 diode
R25732 N25731 N25732 10
D25732 N25732 0 diode
R25733 N25732 N25733 10
D25733 N25733 0 diode
R25734 N25733 N25734 10
D25734 N25734 0 diode
R25735 N25734 N25735 10
D25735 N25735 0 diode
R25736 N25735 N25736 10
D25736 N25736 0 diode
R25737 N25736 N25737 10
D25737 N25737 0 diode
R25738 N25737 N25738 10
D25738 N25738 0 diode
R25739 N25738 N25739 10
D25739 N25739 0 diode
R25740 N25739 N25740 10
D25740 N25740 0 diode
R25741 N25740 N25741 10
D25741 N25741 0 diode
R25742 N25741 N25742 10
D25742 N25742 0 diode
R25743 N25742 N25743 10
D25743 N25743 0 diode
R25744 N25743 N25744 10
D25744 N25744 0 diode
R25745 N25744 N25745 10
D25745 N25745 0 diode
R25746 N25745 N25746 10
D25746 N25746 0 diode
R25747 N25746 N25747 10
D25747 N25747 0 diode
R25748 N25747 N25748 10
D25748 N25748 0 diode
R25749 N25748 N25749 10
D25749 N25749 0 diode
R25750 N25749 N25750 10
D25750 N25750 0 diode
R25751 N25750 N25751 10
D25751 N25751 0 diode
R25752 N25751 N25752 10
D25752 N25752 0 diode
R25753 N25752 N25753 10
D25753 N25753 0 diode
R25754 N25753 N25754 10
D25754 N25754 0 diode
R25755 N25754 N25755 10
D25755 N25755 0 diode
R25756 N25755 N25756 10
D25756 N25756 0 diode
R25757 N25756 N25757 10
D25757 N25757 0 diode
R25758 N25757 N25758 10
D25758 N25758 0 diode
R25759 N25758 N25759 10
D25759 N25759 0 diode
R25760 N25759 N25760 10
D25760 N25760 0 diode
R25761 N25760 N25761 10
D25761 N25761 0 diode
R25762 N25761 N25762 10
D25762 N25762 0 diode
R25763 N25762 N25763 10
D25763 N25763 0 diode
R25764 N25763 N25764 10
D25764 N25764 0 diode
R25765 N25764 N25765 10
D25765 N25765 0 diode
R25766 N25765 N25766 10
D25766 N25766 0 diode
R25767 N25766 N25767 10
D25767 N25767 0 diode
R25768 N25767 N25768 10
D25768 N25768 0 diode
R25769 N25768 N25769 10
D25769 N25769 0 diode
R25770 N25769 N25770 10
D25770 N25770 0 diode
R25771 N25770 N25771 10
D25771 N25771 0 diode
R25772 N25771 N25772 10
D25772 N25772 0 diode
R25773 N25772 N25773 10
D25773 N25773 0 diode
R25774 N25773 N25774 10
D25774 N25774 0 diode
R25775 N25774 N25775 10
D25775 N25775 0 diode
R25776 N25775 N25776 10
D25776 N25776 0 diode
R25777 N25776 N25777 10
D25777 N25777 0 diode
R25778 N25777 N25778 10
D25778 N25778 0 diode
R25779 N25778 N25779 10
D25779 N25779 0 diode
R25780 N25779 N25780 10
D25780 N25780 0 diode
R25781 N25780 N25781 10
D25781 N25781 0 diode
R25782 N25781 N25782 10
D25782 N25782 0 diode
R25783 N25782 N25783 10
D25783 N25783 0 diode
R25784 N25783 N25784 10
D25784 N25784 0 diode
R25785 N25784 N25785 10
D25785 N25785 0 diode
R25786 N25785 N25786 10
D25786 N25786 0 diode
R25787 N25786 N25787 10
D25787 N25787 0 diode
R25788 N25787 N25788 10
D25788 N25788 0 diode
R25789 N25788 N25789 10
D25789 N25789 0 diode
R25790 N25789 N25790 10
D25790 N25790 0 diode
R25791 N25790 N25791 10
D25791 N25791 0 diode
R25792 N25791 N25792 10
D25792 N25792 0 diode
R25793 N25792 N25793 10
D25793 N25793 0 diode
R25794 N25793 N25794 10
D25794 N25794 0 diode
R25795 N25794 N25795 10
D25795 N25795 0 diode
R25796 N25795 N25796 10
D25796 N25796 0 diode
R25797 N25796 N25797 10
D25797 N25797 0 diode
R25798 N25797 N25798 10
D25798 N25798 0 diode
R25799 N25798 N25799 10
D25799 N25799 0 diode
R25800 N25799 N25800 10
D25800 N25800 0 diode
R25801 N25800 N25801 10
D25801 N25801 0 diode
R25802 N25801 N25802 10
D25802 N25802 0 diode
R25803 N25802 N25803 10
D25803 N25803 0 diode
R25804 N25803 N25804 10
D25804 N25804 0 diode
R25805 N25804 N25805 10
D25805 N25805 0 diode
R25806 N25805 N25806 10
D25806 N25806 0 diode
R25807 N25806 N25807 10
D25807 N25807 0 diode
R25808 N25807 N25808 10
D25808 N25808 0 diode
R25809 N25808 N25809 10
D25809 N25809 0 diode
R25810 N25809 N25810 10
D25810 N25810 0 diode
R25811 N25810 N25811 10
D25811 N25811 0 diode
R25812 N25811 N25812 10
D25812 N25812 0 diode
R25813 N25812 N25813 10
D25813 N25813 0 diode
R25814 N25813 N25814 10
D25814 N25814 0 diode
R25815 N25814 N25815 10
D25815 N25815 0 diode
R25816 N25815 N25816 10
D25816 N25816 0 diode
R25817 N25816 N25817 10
D25817 N25817 0 diode
R25818 N25817 N25818 10
D25818 N25818 0 diode
R25819 N25818 N25819 10
D25819 N25819 0 diode
R25820 N25819 N25820 10
D25820 N25820 0 diode
R25821 N25820 N25821 10
D25821 N25821 0 diode
R25822 N25821 N25822 10
D25822 N25822 0 diode
R25823 N25822 N25823 10
D25823 N25823 0 diode
R25824 N25823 N25824 10
D25824 N25824 0 diode
R25825 N25824 N25825 10
D25825 N25825 0 diode
R25826 N25825 N25826 10
D25826 N25826 0 diode
R25827 N25826 N25827 10
D25827 N25827 0 diode
R25828 N25827 N25828 10
D25828 N25828 0 diode
R25829 N25828 N25829 10
D25829 N25829 0 diode
R25830 N25829 N25830 10
D25830 N25830 0 diode
R25831 N25830 N25831 10
D25831 N25831 0 diode
R25832 N25831 N25832 10
D25832 N25832 0 diode
R25833 N25832 N25833 10
D25833 N25833 0 diode
R25834 N25833 N25834 10
D25834 N25834 0 diode
R25835 N25834 N25835 10
D25835 N25835 0 diode
R25836 N25835 N25836 10
D25836 N25836 0 diode
R25837 N25836 N25837 10
D25837 N25837 0 diode
R25838 N25837 N25838 10
D25838 N25838 0 diode
R25839 N25838 N25839 10
D25839 N25839 0 diode
R25840 N25839 N25840 10
D25840 N25840 0 diode
R25841 N25840 N25841 10
D25841 N25841 0 diode
R25842 N25841 N25842 10
D25842 N25842 0 diode
R25843 N25842 N25843 10
D25843 N25843 0 diode
R25844 N25843 N25844 10
D25844 N25844 0 diode
R25845 N25844 N25845 10
D25845 N25845 0 diode
R25846 N25845 N25846 10
D25846 N25846 0 diode
R25847 N25846 N25847 10
D25847 N25847 0 diode
R25848 N25847 N25848 10
D25848 N25848 0 diode
R25849 N25848 N25849 10
D25849 N25849 0 diode
R25850 N25849 N25850 10
D25850 N25850 0 diode
R25851 N25850 N25851 10
D25851 N25851 0 diode
R25852 N25851 N25852 10
D25852 N25852 0 diode
R25853 N25852 N25853 10
D25853 N25853 0 diode
R25854 N25853 N25854 10
D25854 N25854 0 diode
R25855 N25854 N25855 10
D25855 N25855 0 diode
R25856 N25855 N25856 10
D25856 N25856 0 diode
R25857 N25856 N25857 10
D25857 N25857 0 diode
R25858 N25857 N25858 10
D25858 N25858 0 diode
R25859 N25858 N25859 10
D25859 N25859 0 diode
R25860 N25859 N25860 10
D25860 N25860 0 diode
R25861 N25860 N25861 10
D25861 N25861 0 diode
R25862 N25861 N25862 10
D25862 N25862 0 diode
R25863 N25862 N25863 10
D25863 N25863 0 diode
R25864 N25863 N25864 10
D25864 N25864 0 diode
R25865 N25864 N25865 10
D25865 N25865 0 diode
R25866 N25865 N25866 10
D25866 N25866 0 diode
R25867 N25866 N25867 10
D25867 N25867 0 diode
R25868 N25867 N25868 10
D25868 N25868 0 diode
R25869 N25868 N25869 10
D25869 N25869 0 diode
R25870 N25869 N25870 10
D25870 N25870 0 diode
R25871 N25870 N25871 10
D25871 N25871 0 diode
R25872 N25871 N25872 10
D25872 N25872 0 diode
R25873 N25872 N25873 10
D25873 N25873 0 diode
R25874 N25873 N25874 10
D25874 N25874 0 diode
R25875 N25874 N25875 10
D25875 N25875 0 diode
R25876 N25875 N25876 10
D25876 N25876 0 diode
R25877 N25876 N25877 10
D25877 N25877 0 diode
R25878 N25877 N25878 10
D25878 N25878 0 diode
R25879 N25878 N25879 10
D25879 N25879 0 diode
R25880 N25879 N25880 10
D25880 N25880 0 diode
R25881 N25880 N25881 10
D25881 N25881 0 diode
R25882 N25881 N25882 10
D25882 N25882 0 diode
R25883 N25882 N25883 10
D25883 N25883 0 diode
R25884 N25883 N25884 10
D25884 N25884 0 diode
R25885 N25884 N25885 10
D25885 N25885 0 diode
R25886 N25885 N25886 10
D25886 N25886 0 diode
R25887 N25886 N25887 10
D25887 N25887 0 diode
R25888 N25887 N25888 10
D25888 N25888 0 diode
R25889 N25888 N25889 10
D25889 N25889 0 diode
R25890 N25889 N25890 10
D25890 N25890 0 diode
R25891 N25890 N25891 10
D25891 N25891 0 diode
R25892 N25891 N25892 10
D25892 N25892 0 diode
R25893 N25892 N25893 10
D25893 N25893 0 diode
R25894 N25893 N25894 10
D25894 N25894 0 diode
R25895 N25894 N25895 10
D25895 N25895 0 diode
R25896 N25895 N25896 10
D25896 N25896 0 diode
R25897 N25896 N25897 10
D25897 N25897 0 diode
R25898 N25897 N25898 10
D25898 N25898 0 diode
R25899 N25898 N25899 10
D25899 N25899 0 diode
R25900 N25899 N25900 10
D25900 N25900 0 diode
R25901 N25900 N25901 10
D25901 N25901 0 diode
R25902 N25901 N25902 10
D25902 N25902 0 diode
R25903 N25902 N25903 10
D25903 N25903 0 diode
R25904 N25903 N25904 10
D25904 N25904 0 diode
R25905 N25904 N25905 10
D25905 N25905 0 diode
R25906 N25905 N25906 10
D25906 N25906 0 diode
R25907 N25906 N25907 10
D25907 N25907 0 diode
R25908 N25907 N25908 10
D25908 N25908 0 diode
R25909 N25908 N25909 10
D25909 N25909 0 diode
R25910 N25909 N25910 10
D25910 N25910 0 diode
R25911 N25910 N25911 10
D25911 N25911 0 diode
R25912 N25911 N25912 10
D25912 N25912 0 diode
R25913 N25912 N25913 10
D25913 N25913 0 diode
R25914 N25913 N25914 10
D25914 N25914 0 diode
R25915 N25914 N25915 10
D25915 N25915 0 diode
R25916 N25915 N25916 10
D25916 N25916 0 diode
R25917 N25916 N25917 10
D25917 N25917 0 diode
R25918 N25917 N25918 10
D25918 N25918 0 diode
R25919 N25918 N25919 10
D25919 N25919 0 diode
R25920 N25919 N25920 10
D25920 N25920 0 diode
R25921 N25920 N25921 10
D25921 N25921 0 diode
R25922 N25921 N25922 10
D25922 N25922 0 diode
R25923 N25922 N25923 10
D25923 N25923 0 diode
R25924 N25923 N25924 10
D25924 N25924 0 diode
R25925 N25924 N25925 10
D25925 N25925 0 diode
R25926 N25925 N25926 10
D25926 N25926 0 diode
R25927 N25926 N25927 10
D25927 N25927 0 diode
R25928 N25927 N25928 10
D25928 N25928 0 diode
R25929 N25928 N25929 10
D25929 N25929 0 diode
R25930 N25929 N25930 10
D25930 N25930 0 diode
R25931 N25930 N25931 10
D25931 N25931 0 diode
R25932 N25931 N25932 10
D25932 N25932 0 diode
R25933 N25932 N25933 10
D25933 N25933 0 diode
R25934 N25933 N25934 10
D25934 N25934 0 diode
R25935 N25934 N25935 10
D25935 N25935 0 diode
R25936 N25935 N25936 10
D25936 N25936 0 diode
R25937 N25936 N25937 10
D25937 N25937 0 diode
R25938 N25937 N25938 10
D25938 N25938 0 diode
R25939 N25938 N25939 10
D25939 N25939 0 diode
R25940 N25939 N25940 10
D25940 N25940 0 diode
R25941 N25940 N25941 10
D25941 N25941 0 diode
R25942 N25941 N25942 10
D25942 N25942 0 diode
R25943 N25942 N25943 10
D25943 N25943 0 diode
R25944 N25943 N25944 10
D25944 N25944 0 diode
R25945 N25944 N25945 10
D25945 N25945 0 diode
R25946 N25945 N25946 10
D25946 N25946 0 diode
R25947 N25946 N25947 10
D25947 N25947 0 diode
R25948 N25947 N25948 10
D25948 N25948 0 diode
R25949 N25948 N25949 10
D25949 N25949 0 diode
R25950 N25949 N25950 10
D25950 N25950 0 diode
R25951 N25950 N25951 10
D25951 N25951 0 diode
R25952 N25951 N25952 10
D25952 N25952 0 diode
R25953 N25952 N25953 10
D25953 N25953 0 diode
R25954 N25953 N25954 10
D25954 N25954 0 diode
R25955 N25954 N25955 10
D25955 N25955 0 diode
R25956 N25955 N25956 10
D25956 N25956 0 diode
R25957 N25956 N25957 10
D25957 N25957 0 diode
R25958 N25957 N25958 10
D25958 N25958 0 diode
R25959 N25958 N25959 10
D25959 N25959 0 diode
R25960 N25959 N25960 10
D25960 N25960 0 diode
R25961 N25960 N25961 10
D25961 N25961 0 diode
R25962 N25961 N25962 10
D25962 N25962 0 diode
R25963 N25962 N25963 10
D25963 N25963 0 diode
R25964 N25963 N25964 10
D25964 N25964 0 diode
R25965 N25964 N25965 10
D25965 N25965 0 diode
R25966 N25965 N25966 10
D25966 N25966 0 diode
R25967 N25966 N25967 10
D25967 N25967 0 diode
R25968 N25967 N25968 10
D25968 N25968 0 diode
R25969 N25968 N25969 10
D25969 N25969 0 diode
R25970 N25969 N25970 10
D25970 N25970 0 diode
R25971 N25970 N25971 10
D25971 N25971 0 diode
R25972 N25971 N25972 10
D25972 N25972 0 diode
R25973 N25972 N25973 10
D25973 N25973 0 diode
R25974 N25973 N25974 10
D25974 N25974 0 diode
R25975 N25974 N25975 10
D25975 N25975 0 diode
R25976 N25975 N25976 10
D25976 N25976 0 diode
R25977 N25976 N25977 10
D25977 N25977 0 diode
R25978 N25977 N25978 10
D25978 N25978 0 diode
R25979 N25978 N25979 10
D25979 N25979 0 diode
R25980 N25979 N25980 10
D25980 N25980 0 diode
R25981 N25980 N25981 10
D25981 N25981 0 diode
R25982 N25981 N25982 10
D25982 N25982 0 diode
R25983 N25982 N25983 10
D25983 N25983 0 diode
R25984 N25983 N25984 10
D25984 N25984 0 diode
R25985 N25984 N25985 10
D25985 N25985 0 diode
R25986 N25985 N25986 10
D25986 N25986 0 diode
R25987 N25986 N25987 10
D25987 N25987 0 diode
R25988 N25987 N25988 10
D25988 N25988 0 diode
R25989 N25988 N25989 10
D25989 N25989 0 diode
R25990 N25989 N25990 10
D25990 N25990 0 diode
R25991 N25990 N25991 10
D25991 N25991 0 diode
R25992 N25991 N25992 10
D25992 N25992 0 diode
R25993 N25992 N25993 10
D25993 N25993 0 diode
R25994 N25993 N25994 10
D25994 N25994 0 diode
R25995 N25994 N25995 10
D25995 N25995 0 diode
R25996 N25995 N25996 10
D25996 N25996 0 diode
R25997 N25996 N25997 10
D25997 N25997 0 diode
R25998 N25997 N25998 10
D25998 N25998 0 diode
R25999 N25998 N25999 10
D25999 N25999 0 diode
R26000 N25999 N26000 10
D26000 N26000 0 diode
R26001 N26000 N26001 10
D26001 N26001 0 diode
R26002 N26001 N26002 10
D26002 N26002 0 diode
R26003 N26002 N26003 10
D26003 N26003 0 diode
R26004 N26003 N26004 10
D26004 N26004 0 diode
R26005 N26004 N26005 10
D26005 N26005 0 diode
R26006 N26005 N26006 10
D26006 N26006 0 diode
R26007 N26006 N26007 10
D26007 N26007 0 diode
R26008 N26007 N26008 10
D26008 N26008 0 diode
R26009 N26008 N26009 10
D26009 N26009 0 diode
R26010 N26009 N26010 10
D26010 N26010 0 diode
R26011 N26010 N26011 10
D26011 N26011 0 diode
R26012 N26011 N26012 10
D26012 N26012 0 diode
R26013 N26012 N26013 10
D26013 N26013 0 diode
R26014 N26013 N26014 10
D26014 N26014 0 diode
R26015 N26014 N26015 10
D26015 N26015 0 diode
R26016 N26015 N26016 10
D26016 N26016 0 diode
R26017 N26016 N26017 10
D26017 N26017 0 diode
R26018 N26017 N26018 10
D26018 N26018 0 diode
R26019 N26018 N26019 10
D26019 N26019 0 diode
R26020 N26019 N26020 10
D26020 N26020 0 diode
R26021 N26020 N26021 10
D26021 N26021 0 diode
R26022 N26021 N26022 10
D26022 N26022 0 diode
R26023 N26022 N26023 10
D26023 N26023 0 diode
R26024 N26023 N26024 10
D26024 N26024 0 diode
R26025 N26024 N26025 10
D26025 N26025 0 diode
R26026 N26025 N26026 10
D26026 N26026 0 diode
R26027 N26026 N26027 10
D26027 N26027 0 diode
R26028 N26027 N26028 10
D26028 N26028 0 diode
R26029 N26028 N26029 10
D26029 N26029 0 diode
R26030 N26029 N26030 10
D26030 N26030 0 diode
R26031 N26030 N26031 10
D26031 N26031 0 diode
R26032 N26031 N26032 10
D26032 N26032 0 diode
R26033 N26032 N26033 10
D26033 N26033 0 diode
R26034 N26033 N26034 10
D26034 N26034 0 diode
R26035 N26034 N26035 10
D26035 N26035 0 diode
R26036 N26035 N26036 10
D26036 N26036 0 diode
R26037 N26036 N26037 10
D26037 N26037 0 diode
R26038 N26037 N26038 10
D26038 N26038 0 diode
R26039 N26038 N26039 10
D26039 N26039 0 diode
R26040 N26039 N26040 10
D26040 N26040 0 diode
R26041 N26040 N26041 10
D26041 N26041 0 diode
R26042 N26041 N26042 10
D26042 N26042 0 diode
R26043 N26042 N26043 10
D26043 N26043 0 diode
R26044 N26043 N26044 10
D26044 N26044 0 diode
R26045 N26044 N26045 10
D26045 N26045 0 diode
R26046 N26045 N26046 10
D26046 N26046 0 diode
R26047 N26046 N26047 10
D26047 N26047 0 diode
R26048 N26047 N26048 10
D26048 N26048 0 diode
R26049 N26048 N26049 10
D26049 N26049 0 diode
R26050 N26049 N26050 10
D26050 N26050 0 diode
R26051 N26050 N26051 10
D26051 N26051 0 diode
R26052 N26051 N26052 10
D26052 N26052 0 diode
R26053 N26052 N26053 10
D26053 N26053 0 diode
R26054 N26053 N26054 10
D26054 N26054 0 diode
R26055 N26054 N26055 10
D26055 N26055 0 diode
R26056 N26055 N26056 10
D26056 N26056 0 diode
R26057 N26056 N26057 10
D26057 N26057 0 diode
R26058 N26057 N26058 10
D26058 N26058 0 diode
R26059 N26058 N26059 10
D26059 N26059 0 diode
R26060 N26059 N26060 10
D26060 N26060 0 diode
R26061 N26060 N26061 10
D26061 N26061 0 diode
R26062 N26061 N26062 10
D26062 N26062 0 diode
R26063 N26062 N26063 10
D26063 N26063 0 diode
R26064 N26063 N26064 10
D26064 N26064 0 diode
R26065 N26064 N26065 10
D26065 N26065 0 diode
R26066 N26065 N26066 10
D26066 N26066 0 diode
R26067 N26066 N26067 10
D26067 N26067 0 diode
R26068 N26067 N26068 10
D26068 N26068 0 diode
R26069 N26068 N26069 10
D26069 N26069 0 diode
R26070 N26069 N26070 10
D26070 N26070 0 diode
R26071 N26070 N26071 10
D26071 N26071 0 diode
R26072 N26071 N26072 10
D26072 N26072 0 diode
R26073 N26072 N26073 10
D26073 N26073 0 diode
R26074 N26073 N26074 10
D26074 N26074 0 diode
R26075 N26074 N26075 10
D26075 N26075 0 diode
R26076 N26075 N26076 10
D26076 N26076 0 diode
R26077 N26076 N26077 10
D26077 N26077 0 diode
R26078 N26077 N26078 10
D26078 N26078 0 diode
R26079 N26078 N26079 10
D26079 N26079 0 diode
R26080 N26079 N26080 10
D26080 N26080 0 diode
R26081 N26080 N26081 10
D26081 N26081 0 diode
R26082 N26081 N26082 10
D26082 N26082 0 diode
R26083 N26082 N26083 10
D26083 N26083 0 diode
R26084 N26083 N26084 10
D26084 N26084 0 diode
R26085 N26084 N26085 10
D26085 N26085 0 diode
R26086 N26085 N26086 10
D26086 N26086 0 diode
R26087 N26086 N26087 10
D26087 N26087 0 diode
R26088 N26087 N26088 10
D26088 N26088 0 diode
R26089 N26088 N26089 10
D26089 N26089 0 diode
R26090 N26089 N26090 10
D26090 N26090 0 diode
R26091 N26090 N26091 10
D26091 N26091 0 diode
R26092 N26091 N26092 10
D26092 N26092 0 diode
R26093 N26092 N26093 10
D26093 N26093 0 diode
R26094 N26093 N26094 10
D26094 N26094 0 diode
R26095 N26094 N26095 10
D26095 N26095 0 diode
R26096 N26095 N26096 10
D26096 N26096 0 diode
R26097 N26096 N26097 10
D26097 N26097 0 diode
R26098 N26097 N26098 10
D26098 N26098 0 diode
R26099 N26098 N26099 10
D26099 N26099 0 diode
R26100 N26099 N26100 10
D26100 N26100 0 diode
R26101 N26100 N26101 10
D26101 N26101 0 diode
R26102 N26101 N26102 10
D26102 N26102 0 diode
R26103 N26102 N26103 10
D26103 N26103 0 diode
R26104 N26103 N26104 10
D26104 N26104 0 diode
R26105 N26104 N26105 10
D26105 N26105 0 diode
R26106 N26105 N26106 10
D26106 N26106 0 diode
R26107 N26106 N26107 10
D26107 N26107 0 diode
R26108 N26107 N26108 10
D26108 N26108 0 diode
R26109 N26108 N26109 10
D26109 N26109 0 diode
R26110 N26109 N26110 10
D26110 N26110 0 diode
R26111 N26110 N26111 10
D26111 N26111 0 diode
R26112 N26111 N26112 10
D26112 N26112 0 diode
R26113 N26112 N26113 10
D26113 N26113 0 diode
R26114 N26113 N26114 10
D26114 N26114 0 diode
R26115 N26114 N26115 10
D26115 N26115 0 diode
R26116 N26115 N26116 10
D26116 N26116 0 diode
R26117 N26116 N26117 10
D26117 N26117 0 diode
R26118 N26117 N26118 10
D26118 N26118 0 diode
R26119 N26118 N26119 10
D26119 N26119 0 diode
R26120 N26119 N26120 10
D26120 N26120 0 diode
R26121 N26120 N26121 10
D26121 N26121 0 diode
R26122 N26121 N26122 10
D26122 N26122 0 diode
R26123 N26122 N26123 10
D26123 N26123 0 diode
R26124 N26123 N26124 10
D26124 N26124 0 diode
R26125 N26124 N26125 10
D26125 N26125 0 diode
R26126 N26125 N26126 10
D26126 N26126 0 diode
R26127 N26126 N26127 10
D26127 N26127 0 diode
R26128 N26127 N26128 10
D26128 N26128 0 diode
R26129 N26128 N26129 10
D26129 N26129 0 diode
R26130 N26129 N26130 10
D26130 N26130 0 diode
R26131 N26130 N26131 10
D26131 N26131 0 diode
R26132 N26131 N26132 10
D26132 N26132 0 diode
R26133 N26132 N26133 10
D26133 N26133 0 diode
R26134 N26133 N26134 10
D26134 N26134 0 diode
R26135 N26134 N26135 10
D26135 N26135 0 diode
R26136 N26135 N26136 10
D26136 N26136 0 diode
R26137 N26136 N26137 10
D26137 N26137 0 diode
R26138 N26137 N26138 10
D26138 N26138 0 diode
R26139 N26138 N26139 10
D26139 N26139 0 diode
R26140 N26139 N26140 10
D26140 N26140 0 diode
R26141 N26140 N26141 10
D26141 N26141 0 diode
R26142 N26141 N26142 10
D26142 N26142 0 diode
R26143 N26142 N26143 10
D26143 N26143 0 diode
R26144 N26143 N26144 10
D26144 N26144 0 diode
R26145 N26144 N26145 10
D26145 N26145 0 diode
R26146 N26145 N26146 10
D26146 N26146 0 diode
R26147 N26146 N26147 10
D26147 N26147 0 diode
R26148 N26147 N26148 10
D26148 N26148 0 diode
R26149 N26148 N26149 10
D26149 N26149 0 diode
R26150 N26149 N26150 10
D26150 N26150 0 diode
R26151 N26150 N26151 10
D26151 N26151 0 diode
R26152 N26151 N26152 10
D26152 N26152 0 diode
R26153 N26152 N26153 10
D26153 N26153 0 diode
R26154 N26153 N26154 10
D26154 N26154 0 diode
R26155 N26154 N26155 10
D26155 N26155 0 diode
R26156 N26155 N26156 10
D26156 N26156 0 diode
R26157 N26156 N26157 10
D26157 N26157 0 diode
R26158 N26157 N26158 10
D26158 N26158 0 diode
R26159 N26158 N26159 10
D26159 N26159 0 diode
R26160 N26159 N26160 10
D26160 N26160 0 diode
R26161 N26160 N26161 10
D26161 N26161 0 diode
R26162 N26161 N26162 10
D26162 N26162 0 diode
R26163 N26162 N26163 10
D26163 N26163 0 diode
R26164 N26163 N26164 10
D26164 N26164 0 diode
R26165 N26164 N26165 10
D26165 N26165 0 diode
R26166 N26165 N26166 10
D26166 N26166 0 diode
R26167 N26166 N26167 10
D26167 N26167 0 diode
R26168 N26167 N26168 10
D26168 N26168 0 diode
R26169 N26168 N26169 10
D26169 N26169 0 diode
R26170 N26169 N26170 10
D26170 N26170 0 diode
R26171 N26170 N26171 10
D26171 N26171 0 diode
R26172 N26171 N26172 10
D26172 N26172 0 diode
R26173 N26172 N26173 10
D26173 N26173 0 diode
R26174 N26173 N26174 10
D26174 N26174 0 diode
R26175 N26174 N26175 10
D26175 N26175 0 diode
R26176 N26175 N26176 10
D26176 N26176 0 diode
R26177 N26176 N26177 10
D26177 N26177 0 diode
R26178 N26177 N26178 10
D26178 N26178 0 diode
R26179 N26178 N26179 10
D26179 N26179 0 diode
R26180 N26179 N26180 10
D26180 N26180 0 diode
R26181 N26180 N26181 10
D26181 N26181 0 diode
R26182 N26181 N26182 10
D26182 N26182 0 diode
R26183 N26182 N26183 10
D26183 N26183 0 diode
R26184 N26183 N26184 10
D26184 N26184 0 diode
R26185 N26184 N26185 10
D26185 N26185 0 diode
R26186 N26185 N26186 10
D26186 N26186 0 diode
R26187 N26186 N26187 10
D26187 N26187 0 diode
R26188 N26187 N26188 10
D26188 N26188 0 diode
R26189 N26188 N26189 10
D26189 N26189 0 diode
R26190 N26189 N26190 10
D26190 N26190 0 diode
R26191 N26190 N26191 10
D26191 N26191 0 diode
R26192 N26191 N26192 10
D26192 N26192 0 diode
R26193 N26192 N26193 10
D26193 N26193 0 diode
R26194 N26193 N26194 10
D26194 N26194 0 diode
R26195 N26194 N26195 10
D26195 N26195 0 diode
R26196 N26195 N26196 10
D26196 N26196 0 diode
R26197 N26196 N26197 10
D26197 N26197 0 diode
R26198 N26197 N26198 10
D26198 N26198 0 diode
R26199 N26198 N26199 10
D26199 N26199 0 diode
R26200 N26199 N26200 10
D26200 N26200 0 diode
R26201 N26200 N26201 10
D26201 N26201 0 diode
R26202 N26201 N26202 10
D26202 N26202 0 diode
R26203 N26202 N26203 10
D26203 N26203 0 diode
R26204 N26203 N26204 10
D26204 N26204 0 diode
R26205 N26204 N26205 10
D26205 N26205 0 diode
R26206 N26205 N26206 10
D26206 N26206 0 diode
R26207 N26206 N26207 10
D26207 N26207 0 diode
R26208 N26207 N26208 10
D26208 N26208 0 diode
R26209 N26208 N26209 10
D26209 N26209 0 diode
R26210 N26209 N26210 10
D26210 N26210 0 diode
R26211 N26210 N26211 10
D26211 N26211 0 diode
R26212 N26211 N26212 10
D26212 N26212 0 diode
R26213 N26212 N26213 10
D26213 N26213 0 diode
R26214 N26213 N26214 10
D26214 N26214 0 diode
R26215 N26214 N26215 10
D26215 N26215 0 diode
R26216 N26215 N26216 10
D26216 N26216 0 diode
R26217 N26216 N26217 10
D26217 N26217 0 diode
R26218 N26217 N26218 10
D26218 N26218 0 diode
R26219 N26218 N26219 10
D26219 N26219 0 diode
R26220 N26219 N26220 10
D26220 N26220 0 diode
R26221 N26220 N26221 10
D26221 N26221 0 diode
R26222 N26221 N26222 10
D26222 N26222 0 diode
R26223 N26222 N26223 10
D26223 N26223 0 diode
R26224 N26223 N26224 10
D26224 N26224 0 diode
R26225 N26224 N26225 10
D26225 N26225 0 diode
R26226 N26225 N26226 10
D26226 N26226 0 diode
R26227 N26226 N26227 10
D26227 N26227 0 diode
R26228 N26227 N26228 10
D26228 N26228 0 diode
R26229 N26228 N26229 10
D26229 N26229 0 diode
R26230 N26229 N26230 10
D26230 N26230 0 diode
R26231 N26230 N26231 10
D26231 N26231 0 diode
R26232 N26231 N26232 10
D26232 N26232 0 diode
R26233 N26232 N26233 10
D26233 N26233 0 diode
R26234 N26233 N26234 10
D26234 N26234 0 diode
R26235 N26234 N26235 10
D26235 N26235 0 diode
R26236 N26235 N26236 10
D26236 N26236 0 diode
R26237 N26236 N26237 10
D26237 N26237 0 diode
R26238 N26237 N26238 10
D26238 N26238 0 diode
R26239 N26238 N26239 10
D26239 N26239 0 diode
R26240 N26239 N26240 10
D26240 N26240 0 diode
R26241 N26240 N26241 10
D26241 N26241 0 diode
R26242 N26241 N26242 10
D26242 N26242 0 diode
R26243 N26242 N26243 10
D26243 N26243 0 diode
R26244 N26243 N26244 10
D26244 N26244 0 diode
R26245 N26244 N26245 10
D26245 N26245 0 diode
R26246 N26245 N26246 10
D26246 N26246 0 diode
R26247 N26246 N26247 10
D26247 N26247 0 diode
R26248 N26247 N26248 10
D26248 N26248 0 diode
R26249 N26248 N26249 10
D26249 N26249 0 diode
R26250 N26249 N26250 10
D26250 N26250 0 diode
R26251 N26250 N26251 10
D26251 N26251 0 diode
R26252 N26251 N26252 10
D26252 N26252 0 diode
R26253 N26252 N26253 10
D26253 N26253 0 diode
R26254 N26253 N26254 10
D26254 N26254 0 diode
R26255 N26254 N26255 10
D26255 N26255 0 diode
R26256 N26255 N26256 10
D26256 N26256 0 diode
R26257 N26256 N26257 10
D26257 N26257 0 diode
R26258 N26257 N26258 10
D26258 N26258 0 diode
R26259 N26258 N26259 10
D26259 N26259 0 diode
R26260 N26259 N26260 10
D26260 N26260 0 diode
R26261 N26260 N26261 10
D26261 N26261 0 diode
R26262 N26261 N26262 10
D26262 N26262 0 diode
R26263 N26262 N26263 10
D26263 N26263 0 diode
R26264 N26263 N26264 10
D26264 N26264 0 diode
R26265 N26264 N26265 10
D26265 N26265 0 diode
R26266 N26265 N26266 10
D26266 N26266 0 diode
R26267 N26266 N26267 10
D26267 N26267 0 diode
R26268 N26267 N26268 10
D26268 N26268 0 diode
R26269 N26268 N26269 10
D26269 N26269 0 diode
R26270 N26269 N26270 10
D26270 N26270 0 diode
R26271 N26270 N26271 10
D26271 N26271 0 diode
R26272 N26271 N26272 10
D26272 N26272 0 diode
R26273 N26272 N26273 10
D26273 N26273 0 diode
R26274 N26273 N26274 10
D26274 N26274 0 diode
R26275 N26274 N26275 10
D26275 N26275 0 diode
R26276 N26275 N26276 10
D26276 N26276 0 diode
R26277 N26276 N26277 10
D26277 N26277 0 diode
R26278 N26277 N26278 10
D26278 N26278 0 diode
R26279 N26278 N26279 10
D26279 N26279 0 diode
R26280 N26279 N26280 10
D26280 N26280 0 diode
R26281 N26280 N26281 10
D26281 N26281 0 diode
R26282 N26281 N26282 10
D26282 N26282 0 diode
R26283 N26282 N26283 10
D26283 N26283 0 diode
R26284 N26283 N26284 10
D26284 N26284 0 diode
R26285 N26284 N26285 10
D26285 N26285 0 diode
R26286 N26285 N26286 10
D26286 N26286 0 diode
R26287 N26286 N26287 10
D26287 N26287 0 diode
R26288 N26287 N26288 10
D26288 N26288 0 diode
R26289 N26288 N26289 10
D26289 N26289 0 diode
R26290 N26289 N26290 10
D26290 N26290 0 diode
R26291 N26290 N26291 10
D26291 N26291 0 diode
R26292 N26291 N26292 10
D26292 N26292 0 diode
R26293 N26292 N26293 10
D26293 N26293 0 diode
R26294 N26293 N26294 10
D26294 N26294 0 diode
R26295 N26294 N26295 10
D26295 N26295 0 diode
R26296 N26295 N26296 10
D26296 N26296 0 diode
R26297 N26296 N26297 10
D26297 N26297 0 diode
R26298 N26297 N26298 10
D26298 N26298 0 diode
R26299 N26298 N26299 10
D26299 N26299 0 diode
R26300 N26299 N26300 10
D26300 N26300 0 diode
R26301 N26300 N26301 10
D26301 N26301 0 diode
R26302 N26301 N26302 10
D26302 N26302 0 diode
R26303 N26302 N26303 10
D26303 N26303 0 diode
R26304 N26303 N26304 10
D26304 N26304 0 diode
R26305 N26304 N26305 10
D26305 N26305 0 diode
R26306 N26305 N26306 10
D26306 N26306 0 diode
R26307 N26306 N26307 10
D26307 N26307 0 diode
R26308 N26307 N26308 10
D26308 N26308 0 diode
R26309 N26308 N26309 10
D26309 N26309 0 diode
R26310 N26309 N26310 10
D26310 N26310 0 diode
R26311 N26310 N26311 10
D26311 N26311 0 diode
R26312 N26311 N26312 10
D26312 N26312 0 diode
R26313 N26312 N26313 10
D26313 N26313 0 diode
R26314 N26313 N26314 10
D26314 N26314 0 diode
R26315 N26314 N26315 10
D26315 N26315 0 diode
R26316 N26315 N26316 10
D26316 N26316 0 diode
R26317 N26316 N26317 10
D26317 N26317 0 diode
R26318 N26317 N26318 10
D26318 N26318 0 diode
R26319 N26318 N26319 10
D26319 N26319 0 diode
R26320 N26319 N26320 10
D26320 N26320 0 diode
R26321 N26320 N26321 10
D26321 N26321 0 diode
R26322 N26321 N26322 10
D26322 N26322 0 diode
R26323 N26322 N26323 10
D26323 N26323 0 diode
R26324 N26323 N26324 10
D26324 N26324 0 diode
R26325 N26324 N26325 10
D26325 N26325 0 diode
R26326 N26325 N26326 10
D26326 N26326 0 diode
R26327 N26326 N26327 10
D26327 N26327 0 diode
R26328 N26327 N26328 10
D26328 N26328 0 diode
R26329 N26328 N26329 10
D26329 N26329 0 diode
R26330 N26329 N26330 10
D26330 N26330 0 diode
R26331 N26330 N26331 10
D26331 N26331 0 diode
R26332 N26331 N26332 10
D26332 N26332 0 diode
R26333 N26332 N26333 10
D26333 N26333 0 diode
R26334 N26333 N26334 10
D26334 N26334 0 diode
R26335 N26334 N26335 10
D26335 N26335 0 diode
R26336 N26335 N26336 10
D26336 N26336 0 diode
R26337 N26336 N26337 10
D26337 N26337 0 diode
R26338 N26337 N26338 10
D26338 N26338 0 diode
R26339 N26338 N26339 10
D26339 N26339 0 diode
R26340 N26339 N26340 10
D26340 N26340 0 diode
R26341 N26340 N26341 10
D26341 N26341 0 diode
R26342 N26341 N26342 10
D26342 N26342 0 diode
R26343 N26342 N26343 10
D26343 N26343 0 diode
R26344 N26343 N26344 10
D26344 N26344 0 diode
R26345 N26344 N26345 10
D26345 N26345 0 diode
R26346 N26345 N26346 10
D26346 N26346 0 diode
R26347 N26346 N26347 10
D26347 N26347 0 diode
R26348 N26347 N26348 10
D26348 N26348 0 diode
R26349 N26348 N26349 10
D26349 N26349 0 diode
R26350 N26349 N26350 10
D26350 N26350 0 diode
R26351 N26350 N26351 10
D26351 N26351 0 diode
R26352 N26351 N26352 10
D26352 N26352 0 diode
R26353 N26352 N26353 10
D26353 N26353 0 diode
R26354 N26353 N26354 10
D26354 N26354 0 diode
R26355 N26354 N26355 10
D26355 N26355 0 diode
R26356 N26355 N26356 10
D26356 N26356 0 diode
R26357 N26356 N26357 10
D26357 N26357 0 diode
R26358 N26357 N26358 10
D26358 N26358 0 diode
R26359 N26358 N26359 10
D26359 N26359 0 diode
R26360 N26359 N26360 10
D26360 N26360 0 diode
R26361 N26360 N26361 10
D26361 N26361 0 diode
R26362 N26361 N26362 10
D26362 N26362 0 diode
R26363 N26362 N26363 10
D26363 N26363 0 diode
R26364 N26363 N26364 10
D26364 N26364 0 diode
R26365 N26364 N26365 10
D26365 N26365 0 diode
R26366 N26365 N26366 10
D26366 N26366 0 diode
R26367 N26366 N26367 10
D26367 N26367 0 diode
R26368 N26367 N26368 10
D26368 N26368 0 diode
R26369 N26368 N26369 10
D26369 N26369 0 diode
R26370 N26369 N26370 10
D26370 N26370 0 diode
R26371 N26370 N26371 10
D26371 N26371 0 diode
R26372 N26371 N26372 10
D26372 N26372 0 diode
R26373 N26372 N26373 10
D26373 N26373 0 diode
R26374 N26373 N26374 10
D26374 N26374 0 diode
R26375 N26374 N26375 10
D26375 N26375 0 diode
R26376 N26375 N26376 10
D26376 N26376 0 diode
R26377 N26376 N26377 10
D26377 N26377 0 diode
R26378 N26377 N26378 10
D26378 N26378 0 diode
R26379 N26378 N26379 10
D26379 N26379 0 diode
R26380 N26379 N26380 10
D26380 N26380 0 diode
R26381 N26380 N26381 10
D26381 N26381 0 diode
R26382 N26381 N26382 10
D26382 N26382 0 diode
R26383 N26382 N26383 10
D26383 N26383 0 diode
R26384 N26383 N26384 10
D26384 N26384 0 diode
R26385 N26384 N26385 10
D26385 N26385 0 diode
R26386 N26385 N26386 10
D26386 N26386 0 diode
R26387 N26386 N26387 10
D26387 N26387 0 diode
R26388 N26387 N26388 10
D26388 N26388 0 diode
R26389 N26388 N26389 10
D26389 N26389 0 diode
R26390 N26389 N26390 10
D26390 N26390 0 diode
R26391 N26390 N26391 10
D26391 N26391 0 diode
R26392 N26391 N26392 10
D26392 N26392 0 diode
R26393 N26392 N26393 10
D26393 N26393 0 diode
R26394 N26393 N26394 10
D26394 N26394 0 diode
R26395 N26394 N26395 10
D26395 N26395 0 diode
R26396 N26395 N26396 10
D26396 N26396 0 diode
R26397 N26396 N26397 10
D26397 N26397 0 diode
R26398 N26397 N26398 10
D26398 N26398 0 diode
R26399 N26398 N26399 10
D26399 N26399 0 diode
R26400 N26399 N26400 10
D26400 N26400 0 diode
R26401 N26400 N26401 10
D26401 N26401 0 diode
R26402 N26401 N26402 10
D26402 N26402 0 diode
R26403 N26402 N26403 10
D26403 N26403 0 diode
R26404 N26403 N26404 10
D26404 N26404 0 diode
R26405 N26404 N26405 10
D26405 N26405 0 diode
R26406 N26405 N26406 10
D26406 N26406 0 diode
R26407 N26406 N26407 10
D26407 N26407 0 diode
R26408 N26407 N26408 10
D26408 N26408 0 diode
R26409 N26408 N26409 10
D26409 N26409 0 diode
R26410 N26409 N26410 10
D26410 N26410 0 diode
R26411 N26410 N26411 10
D26411 N26411 0 diode
R26412 N26411 N26412 10
D26412 N26412 0 diode
R26413 N26412 N26413 10
D26413 N26413 0 diode
R26414 N26413 N26414 10
D26414 N26414 0 diode
R26415 N26414 N26415 10
D26415 N26415 0 diode
R26416 N26415 N26416 10
D26416 N26416 0 diode
R26417 N26416 N26417 10
D26417 N26417 0 diode
R26418 N26417 N26418 10
D26418 N26418 0 diode
R26419 N26418 N26419 10
D26419 N26419 0 diode
R26420 N26419 N26420 10
D26420 N26420 0 diode
R26421 N26420 N26421 10
D26421 N26421 0 diode
R26422 N26421 N26422 10
D26422 N26422 0 diode
R26423 N26422 N26423 10
D26423 N26423 0 diode
R26424 N26423 N26424 10
D26424 N26424 0 diode
R26425 N26424 N26425 10
D26425 N26425 0 diode
R26426 N26425 N26426 10
D26426 N26426 0 diode
R26427 N26426 N26427 10
D26427 N26427 0 diode
R26428 N26427 N26428 10
D26428 N26428 0 diode
R26429 N26428 N26429 10
D26429 N26429 0 diode
R26430 N26429 N26430 10
D26430 N26430 0 diode
R26431 N26430 N26431 10
D26431 N26431 0 diode
R26432 N26431 N26432 10
D26432 N26432 0 diode
R26433 N26432 N26433 10
D26433 N26433 0 diode
R26434 N26433 N26434 10
D26434 N26434 0 diode
R26435 N26434 N26435 10
D26435 N26435 0 diode
R26436 N26435 N26436 10
D26436 N26436 0 diode
R26437 N26436 N26437 10
D26437 N26437 0 diode
R26438 N26437 N26438 10
D26438 N26438 0 diode
R26439 N26438 N26439 10
D26439 N26439 0 diode
R26440 N26439 N26440 10
D26440 N26440 0 diode
R26441 N26440 N26441 10
D26441 N26441 0 diode
R26442 N26441 N26442 10
D26442 N26442 0 diode
R26443 N26442 N26443 10
D26443 N26443 0 diode
R26444 N26443 N26444 10
D26444 N26444 0 diode
R26445 N26444 N26445 10
D26445 N26445 0 diode
R26446 N26445 N26446 10
D26446 N26446 0 diode
R26447 N26446 N26447 10
D26447 N26447 0 diode
R26448 N26447 N26448 10
D26448 N26448 0 diode
R26449 N26448 N26449 10
D26449 N26449 0 diode
R26450 N26449 N26450 10
D26450 N26450 0 diode
R26451 N26450 N26451 10
D26451 N26451 0 diode
R26452 N26451 N26452 10
D26452 N26452 0 diode
R26453 N26452 N26453 10
D26453 N26453 0 diode
R26454 N26453 N26454 10
D26454 N26454 0 diode
R26455 N26454 N26455 10
D26455 N26455 0 diode
R26456 N26455 N26456 10
D26456 N26456 0 diode
R26457 N26456 N26457 10
D26457 N26457 0 diode
R26458 N26457 N26458 10
D26458 N26458 0 diode
R26459 N26458 N26459 10
D26459 N26459 0 diode
R26460 N26459 N26460 10
D26460 N26460 0 diode
R26461 N26460 N26461 10
D26461 N26461 0 diode
R26462 N26461 N26462 10
D26462 N26462 0 diode
R26463 N26462 N26463 10
D26463 N26463 0 diode
R26464 N26463 N26464 10
D26464 N26464 0 diode
R26465 N26464 N26465 10
D26465 N26465 0 diode
R26466 N26465 N26466 10
D26466 N26466 0 diode
R26467 N26466 N26467 10
D26467 N26467 0 diode
R26468 N26467 N26468 10
D26468 N26468 0 diode
R26469 N26468 N26469 10
D26469 N26469 0 diode
R26470 N26469 N26470 10
D26470 N26470 0 diode
R26471 N26470 N26471 10
D26471 N26471 0 diode
R26472 N26471 N26472 10
D26472 N26472 0 diode
R26473 N26472 N26473 10
D26473 N26473 0 diode
R26474 N26473 N26474 10
D26474 N26474 0 diode
R26475 N26474 N26475 10
D26475 N26475 0 diode
R26476 N26475 N26476 10
D26476 N26476 0 diode
R26477 N26476 N26477 10
D26477 N26477 0 diode
R26478 N26477 N26478 10
D26478 N26478 0 diode
R26479 N26478 N26479 10
D26479 N26479 0 diode
R26480 N26479 N26480 10
D26480 N26480 0 diode
R26481 N26480 N26481 10
D26481 N26481 0 diode
R26482 N26481 N26482 10
D26482 N26482 0 diode
R26483 N26482 N26483 10
D26483 N26483 0 diode
R26484 N26483 N26484 10
D26484 N26484 0 diode
R26485 N26484 N26485 10
D26485 N26485 0 diode
R26486 N26485 N26486 10
D26486 N26486 0 diode
R26487 N26486 N26487 10
D26487 N26487 0 diode
R26488 N26487 N26488 10
D26488 N26488 0 diode
R26489 N26488 N26489 10
D26489 N26489 0 diode
R26490 N26489 N26490 10
D26490 N26490 0 diode
R26491 N26490 N26491 10
D26491 N26491 0 diode
R26492 N26491 N26492 10
D26492 N26492 0 diode
R26493 N26492 N26493 10
D26493 N26493 0 diode
R26494 N26493 N26494 10
D26494 N26494 0 diode
R26495 N26494 N26495 10
D26495 N26495 0 diode
R26496 N26495 N26496 10
D26496 N26496 0 diode
R26497 N26496 N26497 10
D26497 N26497 0 diode
R26498 N26497 N26498 10
D26498 N26498 0 diode
R26499 N26498 N26499 10
D26499 N26499 0 diode
R26500 N26499 N26500 10
D26500 N26500 0 diode
R26501 N26500 N26501 10
D26501 N26501 0 diode
R26502 N26501 N26502 10
D26502 N26502 0 diode
R26503 N26502 N26503 10
D26503 N26503 0 diode
R26504 N26503 N26504 10
D26504 N26504 0 diode
R26505 N26504 N26505 10
D26505 N26505 0 diode
R26506 N26505 N26506 10
D26506 N26506 0 diode
R26507 N26506 N26507 10
D26507 N26507 0 diode
R26508 N26507 N26508 10
D26508 N26508 0 diode
R26509 N26508 N26509 10
D26509 N26509 0 diode
R26510 N26509 N26510 10
D26510 N26510 0 diode
R26511 N26510 N26511 10
D26511 N26511 0 diode
R26512 N26511 N26512 10
D26512 N26512 0 diode
R26513 N26512 N26513 10
D26513 N26513 0 diode
R26514 N26513 N26514 10
D26514 N26514 0 diode
R26515 N26514 N26515 10
D26515 N26515 0 diode
R26516 N26515 N26516 10
D26516 N26516 0 diode
R26517 N26516 N26517 10
D26517 N26517 0 diode
R26518 N26517 N26518 10
D26518 N26518 0 diode
R26519 N26518 N26519 10
D26519 N26519 0 diode
R26520 N26519 N26520 10
D26520 N26520 0 diode
R26521 N26520 N26521 10
D26521 N26521 0 diode
R26522 N26521 N26522 10
D26522 N26522 0 diode
R26523 N26522 N26523 10
D26523 N26523 0 diode
R26524 N26523 N26524 10
D26524 N26524 0 diode
R26525 N26524 N26525 10
D26525 N26525 0 diode
R26526 N26525 N26526 10
D26526 N26526 0 diode
R26527 N26526 N26527 10
D26527 N26527 0 diode
R26528 N26527 N26528 10
D26528 N26528 0 diode
R26529 N26528 N26529 10
D26529 N26529 0 diode
R26530 N26529 N26530 10
D26530 N26530 0 diode
R26531 N26530 N26531 10
D26531 N26531 0 diode
R26532 N26531 N26532 10
D26532 N26532 0 diode
R26533 N26532 N26533 10
D26533 N26533 0 diode
R26534 N26533 N26534 10
D26534 N26534 0 diode
R26535 N26534 N26535 10
D26535 N26535 0 diode
R26536 N26535 N26536 10
D26536 N26536 0 diode
R26537 N26536 N26537 10
D26537 N26537 0 diode
R26538 N26537 N26538 10
D26538 N26538 0 diode
R26539 N26538 N26539 10
D26539 N26539 0 diode
R26540 N26539 N26540 10
D26540 N26540 0 diode
R26541 N26540 N26541 10
D26541 N26541 0 diode
R26542 N26541 N26542 10
D26542 N26542 0 diode
R26543 N26542 N26543 10
D26543 N26543 0 diode
R26544 N26543 N26544 10
D26544 N26544 0 diode
R26545 N26544 N26545 10
D26545 N26545 0 diode
R26546 N26545 N26546 10
D26546 N26546 0 diode
R26547 N26546 N26547 10
D26547 N26547 0 diode
R26548 N26547 N26548 10
D26548 N26548 0 diode
R26549 N26548 N26549 10
D26549 N26549 0 diode
R26550 N26549 N26550 10
D26550 N26550 0 diode
R26551 N26550 N26551 10
D26551 N26551 0 diode
R26552 N26551 N26552 10
D26552 N26552 0 diode
R26553 N26552 N26553 10
D26553 N26553 0 diode
R26554 N26553 N26554 10
D26554 N26554 0 diode
R26555 N26554 N26555 10
D26555 N26555 0 diode
R26556 N26555 N26556 10
D26556 N26556 0 diode
R26557 N26556 N26557 10
D26557 N26557 0 diode
R26558 N26557 N26558 10
D26558 N26558 0 diode
R26559 N26558 N26559 10
D26559 N26559 0 diode
R26560 N26559 N26560 10
D26560 N26560 0 diode
R26561 N26560 N26561 10
D26561 N26561 0 diode
R26562 N26561 N26562 10
D26562 N26562 0 diode
R26563 N26562 N26563 10
D26563 N26563 0 diode
R26564 N26563 N26564 10
D26564 N26564 0 diode
R26565 N26564 N26565 10
D26565 N26565 0 diode
R26566 N26565 N26566 10
D26566 N26566 0 diode
R26567 N26566 N26567 10
D26567 N26567 0 diode
R26568 N26567 N26568 10
D26568 N26568 0 diode
R26569 N26568 N26569 10
D26569 N26569 0 diode
R26570 N26569 N26570 10
D26570 N26570 0 diode
R26571 N26570 N26571 10
D26571 N26571 0 diode
R26572 N26571 N26572 10
D26572 N26572 0 diode
R26573 N26572 N26573 10
D26573 N26573 0 diode
R26574 N26573 N26574 10
D26574 N26574 0 diode
R26575 N26574 N26575 10
D26575 N26575 0 diode
R26576 N26575 N26576 10
D26576 N26576 0 diode
R26577 N26576 N26577 10
D26577 N26577 0 diode
R26578 N26577 N26578 10
D26578 N26578 0 diode
R26579 N26578 N26579 10
D26579 N26579 0 diode
R26580 N26579 N26580 10
D26580 N26580 0 diode
R26581 N26580 N26581 10
D26581 N26581 0 diode
R26582 N26581 N26582 10
D26582 N26582 0 diode
R26583 N26582 N26583 10
D26583 N26583 0 diode
R26584 N26583 N26584 10
D26584 N26584 0 diode
R26585 N26584 N26585 10
D26585 N26585 0 diode
R26586 N26585 N26586 10
D26586 N26586 0 diode
R26587 N26586 N26587 10
D26587 N26587 0 diode
R26588 N26587 N26588 10
D26588 N26588 0 diode
R26589 N26588 N26589 10
D26589 N26589 0 diode
R26590 N26589 N26590 10
D26590 N26590 0 diode
R26591 N26590 N26591 10
D26591 N26591 0 diode
R26592 N26591 N26592 10
D26592 N26592 0 diode
R26593 N26592 N26593 10
D26593 N26593 0 diode
R26594 N26593 N26594 10
D26594 N26594 0 diode
R26595 N26594 N26595 10
D26595 N26595 0 diode
R26596 N26595 N26596 10
D26596 N26596 0 diode
R26597 N26596 N26597 10
D26597 N26597 0 diode
R26598 N26597 N26598 10
D26598 N26598 0 diode
R26599 N26598 N26599 10
D26599 N26599 0 diode
R26600 N26599 N26600 10
D26600 N26600 0 diode
R26601 N26600 N26601 10
D26601 N26601 0 diode
R26602 N26601 N26602 10
D26602 N26602 0 diode
R26603 N26602 N26603 10
D26603 N26603 0 diode
R26604 N26603 N26604 10
D26604 N26604 0 diode
R26605 N26604 N26605 10
D26605 N26605 0 diode
R26606 N26605 N26606 10
D26606 N26606 0 diode
R26607 N26606 N26607 10
D26607 N26607 0 diode
R26608 N26607 N26608 10
D26608 N26608 0 diode
R26609 N26608 N26609 10
D26609 N26609 0 diode
R26610 N26609 N26610 10
D26610 N26610 0 diode
R26611 N26610 N26611 10
D26611 N26611 0 diode
R26612 N26611 N26612 10
D26612 N26612 0 diode
R26613 N26612 N26613 10
D26613 N26613 0 diode
R26614 N26613 N26614 10
D26614 N26614 0 diode
R26615 N26614 N26615 10
D26615 N26615 0 diode
R26616 N26615 N26616 10
D26616 N26616 0 diode
R26617 N26616 N26617 10
D26617 N26617 0 diode
R26618 N26617 N26618 10
D26618 N26618 0 diode
R26619 N26618 N26619 10
D26619 N26619 0 diode
R26620 N26619 N26620 10
D26620 N26620 0 diode
R26621 N26620 N26621 10
D26621 N26621 0 diode
R26622 N26621 N26622 10
D26622 N26622 0 diode
R26623 N26622 N26623 10
D26623 N26623 0 diode
R26624 N26623 N26624 10
D26624 N26624 0 diode
R26625 N26624 N26625 10
D26625 N26625 0 diode
R26626 N26625 N26626 10
D26626 N26626 0 diode
R26627 N26626 N26627 10
D26627 N26627 0 diode
R26628 N26627 N26628 10
D26628 N26628 0 diode
R26629 N26628 N26629 10
D26629 N26629 0 diode
R26630 N26629 N26630 10
D26630 N26630 0 diode
R26631 N26630 N26631 10
D26631 N26631 0 diode
R26632 N26631 N26632 10
D26632 N26632 0 diode
R26633 N26632 N26633 10
D26633 N26633 0 diode
R26634 N26633 N26634 10
D26634 N26634 0 diode
R26635 N26634 N26635 10
D26635 N26635 0 diode
R26636 N26635 N26636 10
D26636 N26636 0 diode
R26637 N26636 N26637 10
D26637 N26637 0 diode
R26638 N26637 N26638 10
D26638 N26638 0 diode
R26639 N26638 N26639 10
D26639 N26639 0 diode
R26640 N26639 N26640 10
D26640 N26640 0 diode
R26641 N26640 N26641 10
D26641 N26641 0 diode
R26642 N26641 N26642 10
D26642 N26642 0 diode
R26643 N26642 N26643 10
D26643 N26643 0 diode
R26644 N26643 N26644 10
D26644 N26644 0 diode
R26645 N26644 N26645 10
D26645 N26645 0 diode
R26646 N26645 N26646 10
D26646 N26646 0 diode
R26647 N26646 N26647 10
D26647 N26647 0 diode
R26648 N26647 N26648 10
D26648 N26648 0 diode
R26649 N26648 N26649 10
D26649 N26649 0 diode
R26650 N26649 N26650 10
D26650 N26650 0 diode
R26651 N26650 N26651 10
D26651 N26651 0 diode
R26652 N26651 N26652 10
D26652 N26652 0 diode
R26653 N26652 N26653 10
D26653 N26653 0 diode
R26654 N26653 N26654 10
D26654 N26654 0 diode
R26655 N26654 N26655 10
D26655 N26655 0 diode
R26656 N26655 N26656 10
D26656 N26656 0 diode
R26657 N26656 N26657 10
D26657 N26657 0 diode
R26658 N26657 N26658 10
D26658 N26658 0 diode
R26659 N26658 N26659 10
D26659 N26659 0 diode
R26660 N26659 N26660 10
D26660 N26660 0 diode
R26661 N26660 N26661 10
D26661 N26661 0 diode
R26662 N26661 N26662 10
D26662 N26662 0 diode
R26663 N26662 N26663 10
D26663 N26663 0 diode
R26664 N26663 N26664 10
D26664 N26664 0 diode
R26665 N26664 N26665 10
D26665 N26665 0 diode
R26666 N26665 N26666 10
D26666 N26666 0 diode
R26667 N26666 N26667 10
D26667 N26667 0 diode
R26668 N26667 N26668 10
D26668 N26668 0 diode
R26669 N26668 N26669 10
D26669 N26669 0 diode
R26670 N26669 N26670 10
D26670 N26670 0 diode
R26671 N26670 N26671 10
D26671 N26671 0 diode
R26672 N26671 N26672 10
D26672 N26672 0 diode
R26673 N26672 N26673 10
D26673 N26673 0 diode
R26674 N26673 N26674 10
D26674 N26674 0 diode
R26675 N26674 N26675 10
D26675 N26675 0 diode
R26676 N26675 N26676 10
D26676 N26676 0 diode
R26677 N26676 N26677 10
D26677 N26677 0 diode
R26678 N26677 N26678 10
D26678 N26678 0 diode
R26679 N26678 N26679 10
D26679 N26679 0 diode
R26680 N26679 N26680 10
D26680 N26680 0 diode
R26681 N26680 N26681 10
D26681 N26681 0 diode
R26682 N26681 N26682 10
D26682 N26682 0 diode
R26683 N26682 N26683 10
D26683 N26683 0 diode
R26684 N26683 N26684 10
D26684 N26684 0 diode
R26685 N26684 N26685 10
D26685 N26685 0 diode
R26686 N26685 N26686 10
D26686 N26686 0 diode
R26687 N26686 N26687 10
D26687 N26687 0 diode
R26688 N26687 N26688 10
D26688 N26688 0 diode
R26689 N26688 N26689 10
D26689 N26689 0 diode
R26690 N26689 N26690 10
D26690 N26690 0 diode
R26691 N26690 N26691 10
D26691 N26691 0 diode
R26692 N26691 N26692 10
D26692 N26692 0 diode
R26693 N26692 N26693 10
D26693 N26693 0 diode
R26694 N26693 N26694 10
D26694 N26694 0 diode
R26695 N26694 N26695 10
D26695 N26695 0 diode
R26696 N26695 N26696 10
D26696 N26696 0 diode
R26697 N26696 N26697 10
D26697 N26697 0 diode
R26698 N26697 N26698 10
D26698 N26698 0 diode
R26699 N26698 N26699 10
D26699 N26699 0 diode
R26700 N26699 N26700 10
D26700 N26700 0 diode
R26701 N26700 N26701 10
D26701 N26701 0 diode
R26702 N26701 N26702 10
D26702 N26702 0 diode
R26703 N26702 N26703 10
D26703 N26703 0 diode
R26704 N26703 N26704 10
D26704 N26704 0 diode
R26705 N26704 N26705 10
D26705 N26705 0 diode
R26706 N26705 N26706 10
D26706 N26706 0 diode
R26707 N26706 N26707 10
D26707 N26707 0 diode
R26708 N26707 N26708 10
D26708 N26708 0 diode
R26709 N26708 N26709 10
D26709 N26709 0 diode
R26710 N26709 N26710 10
D26710 N26710 0 diode
R26711 N26710 N26711 10
D26711 N26711 0 diode
R26712 N26711 N26712 10
D26712 N26712 0 diode
R26713 N26712 N26713 10
D26713 N26713 0 diode
R26714 N26713 N26714 10
D26714 N26714 0 diode
R26715 N26714 N26715 10
D26715 N26715 0 diode
R26716 N26715 N26716 10
D26716 N26716 0 diode
R26717 N26716 N26717 10
D26717 N26717 0 diode
R26718 N26717 N26718 10
D26718 N26718 0 diode
R26719 N26718 N26719 10
D26719 N26719 0 diode
R26720 N26719 N26720 10
D26720 N26720 0 diode
R26721 N26720 N26721 10
D26721 N26721 0 diode
R26722 N26721 N26722 10
D26722 N26722 0 diode
R26723 N26722 N26723 10
D26723 N26723 0 diode
R26724 N26723 N26724 10
D26724 N26724 0 diode
R26725 N26724 N26725 10
D26725 N26725 0 diode
R26726 N26725 N26726 10
D26726 N26726 0 diode
R26727 N26726 N26727 10
D26727 N26727 0 diode
R26728 N26727 N26728 10
D26728 N26728 0 diode
R26729 N26728 N26729 10
D26729 N26729 0 diode
R26730 N26729 N26730 10
D26730 N26730 0 diode
R26731 N26730 N26731 10
D26731 N26731 0 diode
R26732 N26731 N26732 10
D26732 N26732 0 diode
R26733 N26732 N26733 10
D26733 N26733 0 diode
R26734 N26733 N26734 10
D26734 N26734 0 diode
R26735 N26734 N26735 10
D26735 N26735 0 diode
R26736 N26735 N26736 10
D26736 N26736 0 diode
R26737 N26736 N26737 10
D26737 N26737 0 diode
R26738 N26737 N26738 10
D26738 N26738 0 diode
R26739 N26738 N26739 10
D26739 N26739 0 diode
R26740 N26739 N26740 10
D26740 N26740 0 diode
R26741 N26740 N26741 10
D26741 N26741 0 diode
R26742 N26741 N26742 10
D26742 N26742 0 diode
R26743 N26742 N26743 10
D26743 N26743 0 diode
R26744 N26743 N26744 10
D26744 N26744 0 diode
R26745 N26744 N26745 10
D26745 N26745 0 diode
R26746 N26745 N26746 10
D26746 N26746 0 diode
R26747 N26746 N26747 10
D26747 N26747 0 diode
R26748 N26747 N26748 10
D26748 N26748 0 diode
R26749 N26748 N26749 10
D26749 N26749 0 diode
R26750 N26749 N26750 10
D26750 N26750 0 diode
R26751 N26750 N26751 10
D26751 N26751 0 diode
R26752 N26751 N26752 10
D26752 N26752 0 diode
R26753 N26752 N26753 10
D26753 N26753 0 diode
R26754 N26753 N26754 10
D26754 N26754 0 diode
R26755 N26754 N26755 10
D26755 N26755 0 diode
R26756 N26755 N26756 10
D26756 N26756 0 diode
R26757 N26756 N26757 10
D26757 N26757 0 diode
R26758 N26757 N26758 10
D26758 N26758 0 diode
R26759 N26758 N26759 10
D26759 N26759 0 diode
R26760 N26759 N26760 10
D26760 N26760 0 diode
R26761 N26760 N26761 10
D26761 N26761 0 diode
R26762 N26761 N26762 10
D26762 N26762 0 diode
R26763 N26762 N26763 10
D26763 N26763 0 diode
R26764 N26763 N26764 10
D26764 N26764 0 diode
R26765 N26764 N26765 10
D26765 N26765 0 diode
R26766 N26765 N26766 10
D26766 N26766 0 diode
R26767 N26766 N26767 10
D26767 N26767 0 diode
R26768 N26767 N26768 10
D26768 N26768 0 diode
R26769 N26768 N26769 10
D26769 N26769 0 diode
R26770 N26769 N26770 10
D26770 N26770 0 diode
R26771 N26770 N26771 10
D26771 N26771 0 diode
R26772 N26771 N26772 10
D26772 N26772 0 diode
R26773 N26772 N26773 10
D26773 N26773 0 diode
R26774 N26773 N26774 10
D26774 N26774 0 diode
R26775 N26774 N26775 10
D26775 N26775 0 diode
R26776 N26775 N26776 10
D26776 N26776 0 diode
R26777 N26776 N26777 10
D26777 N26777 0 diode
R26778 N26777 N26778 10
D26778 N26778 0 diode
R26779 N26778 N26779 10
D26779 N26779 0 diode
R26780 N26779 N26780 10
D26780 N26780 0 diode
R26781 N26780 N26781 10
D26781 N26781 0 diode
R26782 N26781 N26782 10
D26782 N26782 0 diode
R26783 N26782 N26783 10
D26783 N26783 0 diode
R26784 N26783 N26784 10
D26784 N26784 0 diode
R26785 N26784 N26785 10
D26785 N26785 0 diode
R26786 N26785 N26786 10
D26786 N26786 0 diode
R26787 N26786 N26787 10
D26787 N26787 0 diode
R26788 N26787 N26788 10
D26788 N26788 0 diode
R26789 N26788 N26789 10
D26789 N26789 0 diode
R26790 N26789 N26790 10
D26790 N26790 0 diode
R26791 N26790 N26791 10
D26791 N26791 0 diode
R26792 N26791 N26792 10
D26792 N26792 0 diode
R26793 N26792 N26793 10
D26793 N26793 0 diode
R26794 N26793 N26794 10
D26794 N26794 0 diode
R26795 N26794 N26795 10
D26795 N26795 0 diode
R26796 N26795 N26796 10
D26796 N26796 0 diode
R26797 N26796 N26797 10
D26797 N26797 0 diode
R26798 N26797 N26798 10
D26798 N26798 0 diode
R26799 N26798 N26799 10
D26799 N26799 0 diode
R26800 N26799 N26800 10
D26800 N26800 0 diode
R26801 N26800 N26801 10
D26801 N26801 0 diode
R26802 N26801 N26802 10
D26802 N26802 0 diode
R26803 N26802 N26803 10
D26803 N26803 0 diode
R26804 N26803 N26804 10
D26804 N26804 0 diode
R26805 N26804 N26805 10
D26805 N26805 0 diode
R26806 N26805 N26806 10
D26806 N26806 0 diode
R26807 N26806 N26807 10
D26807 N26807 0 diode
R26808 N26807 N26808 10
D26808 N26808 0 diode
R26809 N26808 N26809 10
D26809 N26809 0 diode
R26810 N26809 N26810 10
D26810 N26810 0 diode
R26811 N26810 N26811 10
D26811 N26811 0 diode
R26812 N26811 N26812 10
D26812 N26812 0 diode
R26813 N26812 N26813 10
D26813 N26813 0 diode
R26814 N26813 N26814 10
D26814 N26814 0 diode
R26815 N26814 N26815 10
D26815 N26815 0 diode
R26816 N26815 N26816 10
D26816 N26816 0 diode
R26817 N26816 N26817 10
D26817 N26817 0 diode
R26818 N26817 N26818 10
D26818 N26818 0 diode
R26819 N26818 N26819 10
D26819 N26819 0 diode
R26820 N26819 N26820 10
D26820 N26820 0 diode
R26821 N26820 N26821 10
D26821 N26821 0 diode
R26822 N26821 N26822 10
D26822 N26822 0 diode
R26823 N26822 N26823 10
D26823 N26823 0 diode
R26824 N26823 N26824 10
D26824 N26824 0 diode
R26825 N26824 N26825 10
D26825 N26825 0 diode
R26826 N26825 N26826 10
D26826 N26826 0 diode
R26827 N26826 N26827 10
D26827 N26827 0 diode
R26828 N26827 N26828 10
D26828 N26828 0 diode
R26829 N26828 N26829 10
D26829 N26829 0 diode
R26830 N26829 N26830 10
D26830 N26830 0 diode
R26831 N26830 N26831 10
D26831 N26831 0 diode
R26832 N26831 N26832 10
D26832 N26832 0 diode
R26833 N26832 N26833 10
D26833 N26833 0 diode
R26834 N26833 N26834 10
D26834 N26834 0 diode
R26835 N26834 N26835 10
D26835 N26835 0 diode
R26836 N26835 N26836 10
D26836 N26836 0 diode
R26837 N26836 N26837 10
D26837 N26837 0 diode
R26838 N26837 N26838 10
D26838 N26838 0 diode
R26839 N26838 N26839 10
D26839 N26839 0 diode
R26840 N26839 N26840 10
D26840 N26840 0 diode
R26841 N26840 N26841 10
D26841 N26841 0 diode
R26842 N26841 N26842 10
D26842 N26842 0 diode
R26843 N26842 N26843 10
D26843 N26843 0 diode
R26844 N26843 N26844 10
D26844 N26844 0 diode
R26845 N26844 N26845 10
D26845 N26845 0 diode
R26846 N26845 N26846 10
D26846 N26846 0 diode
R26847 N26846 N26847 10
D26847 N26847 0 diode
R26848 N26847 N26848 10
D26848 N26848 0 diode
R26849 N26848 N26849 10
D26849 N26849 0 diode
R26850 N26849 N26850 10
D26850 N26850 0 diode
R26851 N26850 N26851 10
D26851 N26851 0 diode
R26852 N26851 N26852 10
D26852 N26852 0 diode
R26853 N26852 N26853 10
D26853 N26853 0 diode
R26854 N26853 N26854 10
D26854 N26854 0 diode
R26855 N26854 N26855 10
D26855 N26855 0 diode
R26856 N26855 N26856 10
D26856 N26856 0 diode
R26857 N26856 N26857 10
D26857 N26857 0 diode
R26858 N26857 N26858 10
D26858 N26858 0 diode
R26859 N26858 N26859 10
D26859 N26859 0 diode
R26860 N26859 N26860 10
D26860 N26860 0 diode
R26861 N26860 N26861 10
D26861 N26861 0 diode
R26862 N26861 N26862 10
D26862 N26862 0 diode
R26863 N26862 N26863 10
D26863 N26863 0 diode
R26864 N26863 N26864 10
D26864 N26864 0 diode
R26865 N26864 N26865 10
D26865 N26865 0 diode
R26866 N26865 N26866 10
D26866 N26866 0 diode
R26867 N26866 N26867 10
D26867 N26867 0 diode
R26868 N26867 N26868 10
D26868 N26868 0 diode
R26869 N26868 N26869 10
D26869 N26869 0 diode
R26870 N26869 N26870 10
D26870 N26870 0 diode
R26871 N26870 N26871 10
D26871 N26871 0 diode
R26872 N26871 N26872 10
D26872 N26872 0 diode
R26873 N26872 N26873 10
D26873 N26873 0 diode
R26874 N26873 N26874 10
D26874 N26874 0 diode
R26875 N26874 N26875 10
D26875 N26875 0 diode
R26876 N26875 N26876 10
D26876 N26876 0 diode
R26877 N26876 N26877 10
D26877 N26877 0 diode
R26878 N26877 N26878 10
D26878 N26878 0 diode
R26879 N26878 N26879 10
D26879 N26879 0 diode
R26880 N26879 N26880 10
D26880 N26880 0 diode
R26881 N26880 N26881 10
D26881 N26881 0 diode
R26882 N26881 N26882 10
D26882 N26882 0 diode
R26883 N26882 N26883 10
D26883 N26883 0 diode
R26884 N26883 N26884 10
D26884 N26884 0 diode
R26885 N26884 N26885 10
D26885 N26885 0 diode
R26886 N26885 N26886 10
D26886 N26886 0 diode
R26887 N26886 N26887 10
D26887 N26887 0 diode
R26888 N26887 N26888 10
D26888 N26888 0 diode
R26889 N26888 N26889 10
D26889 N26889 0 diode
R26890 N26889 N26890 10
D26890 N26890 0 diode
R26891 N26890 N26891 10
D26891 N26891 0 diode
R26892 N26891 N26892 10
D26892 N26892 0 diode
R26893 N26892 N26893 10
D26893 N26893 0 diode
R26894 N26893 N26894 10
D26894 N26894 0 diode
R26895 N26894 N26895 10
D26895 N26895 0 diode
R26896 N26895 N26896 10
D26896 N26896 0 diode
R26897 N26896 N26897 10
D26897 N26897 0 diode
R26898 N26897 N26898 10
D26898 N26898 0 diode
R26899 N26898 N26899 10
D26899 N26899 0 diode
R26900 N26899 N26900 10
D26900 N26900 0 diode
R26901 N26900 N26901 10
D26901 N26901 0 diode
R26902 N26901 N26902 10
D26902 N26902 0 diode
R26903 N26902 N26903 10
D26903 N26903 0 diode
R26904 N26903 N26904 10
D26904 N26904 0 diode
R26905 N26904 N26905 10
D26905 N26905 0 diode
R26906 N26905 N26906 10
D26906 N26906 0 diode
R26907 N26906 N26907 10
D26907 N26907 0 diode
R26908 N26907 N26908 10
D26908 N26908 0 diode
R26909 N26908 N26909 10
D26909 N26909 0 diode
R26910 N26909 N26910 10
D26910 N26910 0 diode
R26911 N26910 N26911 10
D26911 N26911 0 diode
R26912 N26911 N26912 10
D26912 N26912 0 diode
R26913 N26912 N26913 10
D26913 N26913 0 diode
R26914 N26913 N26914 10
D26914 N26914 0 diode
R26915 N26914 N26915 10
D26915 N26915 0 diode
R26916 N26915 N26916 10
D26916 N26916 0 diode
R26917 N26916 N26917 10
D26917 N26917 0 diode
R26918 N26917 N26918 10
D26918 N26918 0 diode
R26919 N26918 N26919 10
D26919 N26919 0 diode
R26920 N26919 N26920 10
D26920 N26920 0 diode
R26921 N26920 N26921 10
D26921 N26921 0 diode
R26922 N26921 N26922 10
D26922 N26922 0 diode
R26923 N26922 N26923 10
D26923 N26923 0 diode
R26924 N26923 N26924 10
D26924 N26924 0 diode
R26925 N26924 N26925 10
D26925 N26925 0 diode
R26926 N26925 N26926 10
D26926 N26926 0 diode
R26927 N26926 N26927 10
D26927 N26927 0 diode
R26928 N26927 N26928 10
D26928 N26928 0 diode
R26929 N26928 N26929 10
D26929 N26929 0 diode
R26930 N26929 N26930 10
D26930 N26930 0 diode
R26931 N26930 N26931 10
D26931 N26931 0 diode
R26932 N26931 N26932 10
D26932 N26932 0 diode
R26933 N26932 N26933 10
D26933 N26933 0 diode
R26934 N26933 N26934 10
D26934 N26934 0 diode
R26935 N26934 N26935 10
D26935 N26935 0 diode
R26936 N26935 N26936 10
D26936 N26936 0 diode
R26937 N26936 N26937 10
D26937 N26937 0 diode
R26938 N26937 N26938 10
D26938 N26938 0 diode
R26939 N26938 N26939 10
D26939 N26939 0 diode
R26940 N26939 N26940 10
D26940 N26940 0 diode
R26941 N26940 N26941 10
D26941 N26941 0 diode
R26942 N26941 N26942 10
D26942 N26942 0 diode
R26943 N26942 N26943 10
D26943 N26943 0 diode
R26944 N26943 N26944 10
D26944 N26944 0 diode
R26945 N26944 N26945 10
D26945 N26945 0 diode
R26946 N26945 N26946 10
D26946 N26946 0 diode
R26947 N26946 N26947 10
D26947 N26947 0 diode
R26948 N26947 N26948 10
D26948 N26948 0 diode
R26949 N26948 N26949 10
D26949 N26949 0 diode
R26950 N26949 N26950 10
D26950 N26950 0 diode
R26951 N26950 N26951 10
D26951 N26951 0 diode
R26952 N26951 N26952 10
D26952 N26952 0 diode
R26953 N26952 N26953 10
D26953 N26953 0 diode
R26954 N26953 N26954 10
D26954 N26954 0 diode
R26955 N26954 N26955 10
D26955 N26955 0 diode
R26956 N26955 N26956 10
D26956 N26956 0 diode
R26957 N26956 N26957 10
D26957 N26957 0 diode
R26958 N26957 N26958 10
D26958 N26958 0 diode
R26959 N26958 N26959 10
D26959 N26959 0 diode
R26960 N26959 N26960 10
D26960 N26960 0 diode
R26961 N26960 N26961 10
D26961 N26961 0 diode
R26962 N26961 N26962 10
D26962 N26962 0 diode
R26963 N26962 N26963 10
D26963 N26963 0 diode
R26964 N26963 N26964 10
D26964 N26964 0 diode
R26965 N26964 N26965 10
D26965 N26965 0 diode
R26966 N26965 N26966 10
D26966 N26966 0 diode
R26967 N26966 N26967 10
D26967 N26967 0 diode
R26968 N26967 N26968 10
D26968 N26968 0 diode
R26969 N26968 N26969 10
D26969 N26969 0 diode
R26970 N26969 N26970 10
D26970 N26970 0 diode
R26971 N26970 N26971 10
D26971 N26971 0 diode
R26972 N26971 N26972 10
D26972 N26972 0 diode
R26973 N26972 N26973 10
D26973 N26973 0 diode
R26974 N26973 N26974 10
D26974 N26974 0 diode
R26975 N26974 N26975 10
D26975 N26975 0 diode
R26976 N26975 N26976 10
D26976 N26976 0 diode
R26977 N26976 N26977 10
D26977 N26977 0 diode
R26978 N26977 N26978 10
D26978 N26978 0 diode
R26979 N26978 N26979 10
D26979 N26979 0 diode
R26980 N26979 N26980 10
D26980 N26980 0 diode
R26981 N26980 N26981 10
D26981 N26981 0 diode
R26982 N26981 N26982 10
D26982 N26982 0 diode
R26983 N26982 N26983 10
D26983 N26983 0 diode
R26984 N26983 N26984 10
D26984 N26984 0 diode
R26985 N26984 N26985 10
D26985 N26985 0 diode
R26986 N26985 N26986 10
D26986 N26986 0 diode
R26987 N26986 N26987 10
D26987 N26987 0 diode
R26988 N26987 N26988 10
D26988 N26988 0 diode
R26989 N26988 N26989 10
D26989 N26989 0 diode
R26990 N26989 N26990 10
D26990 N26990 0 diode
R26991 N26990 N26991 10
D26991 N26991 0 diode
R26992 N26991 N26992 10
D26992 N26992 0 diode
R26993 N26992 N26993 10
D26993 N26993 0 diode
R26994 N26993 N26994 10
D26994 N26994 0 diode
R26995 N26994 N26995 10
D26995 N26995 0 diode
R26996 N26995 N26996 10
D26996 N26996 0 diode
R26997 N26996 N26997 10
D26997 N26997 0 diode
R26998 N26997 N26998 10
D26998 N26998 0 diode
R26999 N26998 N26999 10
D26999 N26999 0 diode
R27000 N26999 N27000 10
D27000 N27000 0 diode
R27001 N27000 N27001 10
D27001 N27001 0 diode
R27002 N27001 N27002 10
D27002 N27002 0 diode
R27003 N27002 N27003 10
D27003 N27003 0 diode
R27004 N27003 N27004 10
D27004 N27004 0 diode
R27005 N27004 N27005 10
D27005 N27005 0 diode
R27006 N27005 N27006 10
D27006 N27006 0 diode
R27007 N27006 N27007 10
D27007 N27007 0 diode
R27008 N27007 N27008 10
D27008 N27008 0 diode
R27009 N27008 N27009 10
D27009 N27009 0 diode
R27010 N27009 N27010 10
D27010 N27010 0 diode
R27011 N27010 N27011 10
D27011 N27011 0 diode
R27012 N27011 N27012 10
D27012 N27012 0 diode
R27013 N27012 N27013 10
D27013 N27013 0 diode
R27014 N27013 N27014 10
D27014 N27014 0 diode
R27015 N27014 N27015 10
D27015 N27015 0 diode
R27016 N27015 N27016 10
D27016 N27016 0 diode
R27017 N27016 N27017 10
D27017 N27017 0 diode
R27018 N27017 N27018 10
D27018 N27018 0 diode
R27019 N27018 N27019 10
D27019 N27019 0 diode
R27020 N27019 N27020 10
D27020 N27020 0 diode
R27021 N27020 N27021 10
D27021 N27021 0 diode
R27022 N27021 N27022 10
D27022 N27022 0 diode
R27023 N27022 N27023 10
D27023 N27023 0 diode
R27024 N27023 N27024 10
D27024 N27024 0 diode
R27025 N27024 N27025 10
D27025 N27025 0 diode
R27026 N27025 N27026 10
D27026 N27026 0 diode
R27027 N27026 N27027 10
D27027 N27027 0 diode
R27028 N27027 N27028 10
D27028 N27028 0 diode
R27029 N27028 N27029 10
D27029 N27029 0 diode
R27030 N27029 N27030 10
D27030 N27030 0 diode
R27031 N27030 N27031 10
D27031 N27031 0 diode
R27032 N27031 N27032 10
D27032 N27032 0 diode
R27033 N27032 N27033 10
D27033 N27033 0 diode
R27034 N27033 N27034 10
D27034 N27034 0 diode
R27035 N27034 N27035 10
D27035 N27035 0 diode
R27036 N27035 N27036 10
D27036 N27036 0 diode
R27037 N27036 N27037 10
D27037 N27037 0 diode
R27038 N27037 N27038 10
D27038 N27038 0 diode
R27039 N27038 N27039 10
D27039 N27039 0 diode
R27040 N27039 N27040 10
D27040 N27040 0 diode
R27041 N27040 N27041 10
D27041 N27041 0 diode
R27042 N27041 N27042 10
D27042 N27042 0 diode
R27043 N27042 N27043 10
D27043 N27043 0 diode
R27044 N27043 N27044 10
D27044 N27044 0 diode
R27045 N27044 N27045 10
D27045 N27045 0 diode
R27046 N27045 N27046 10
D27046 N27046 0 diode
R27047 N27046 N27047 10
D27047 N27047 0 diode
R27048 N27047 N27048 10
D27048 N27048 0 diode
R27049 N27048 N27049 10
D27049 N27049 0 diode
R27050 N27049 N27050 10
D27050 N27050 0 diode
R27051 N27050 N27051 10
D27051 N27051 0 diode
R27052 N27051 N27052 10
D27052 N27052 0 diode
R27053 N27052 N27053 10
D27053 N27053 0 diode
R27054 N27053 N27054 10
D27054 N27054 0 diode
R27055 N27054 N27055 10
D27055 N27055 0 diode
R27056 N27055 N27056 10
D27056 N27056 0 diode
R27057 N27056 N27057 10
D27057 N27057 0 diode
R27058 N27057 N27058 10
D27058 N27058 0 diode
R27059 N27058 N27059 10
D27059 N27059 0 diode
R27060 N27059 N27060 10
D27060 N27060 0 diode
R27061 N27060 N27061 10
D27061 N27061 0 diode
R27062 N27061 N27062 10
D27062 N27062 0 diode
R27063 N27062 N27063 10
D27063 N27063 0 diode
R27064 N27063 N27064 10
D27064 N27064 0 diode
R27065 N27064 N27065 10
D27065 N27065 0 diode
R27066 N27065 N27066 10
D27066 N27066 0 diode
R27067 N27066 N27067 10
D27067 N27067 0 diode
R27068 N27067 N27068 10
D27068 N27068 0 diode
R27069 N27068 N27069 10
D27069 N27069 0 diode
R27070 N27069 N27070 10
D27070 N27070 0 diode
R27071 N27070 N27071 10
D27071 N27071 0 diode
R27072 N27071 N27072 10
D27072 N27072 0 diode
R27073 N27072 N27073 10
D27073 N27073 0 diode
R27074 N27073 N27074 10
D27074 N27074 0 diode
R27075 N27074 N27075 10
D27075 N27075 0 diode
R27076 N27075 N27076 10
D27076 N27076 0 diode
R27077 N27076 N27077 10
D27077 N27077 0 diode
R27078 N27077 N27078 10
D27078 N27078 0 diode
R27079 N27078 N27079 10
D27079 N27079 0 diode
R27080 N27079 N27080 10
D27080 N27080 0 diode
R27081 N27080 N27081 10
D27081 N27081 0 diode
R27082 N27081 N27082 10
D27082 N27082 0 diode
R27083 N27082 N27083 10
D27083 N27083 0 diode
R27084 N27083 N27084 10
D27084 N27084 0 diode
R27085 N27084 N27085 10
D27085 N27085 0 diode
R27086 N27085 N27086 10
D27086 N27086 0 diode
R27087 N27086 N27087 10
D27087 N27087 0 diode
R27088 N27087 N27088 10
D27088 N27088 0 diode
R27089 N27088 N27089 10
D27089 N27089 0 diode
R27090 N27089 N27090 10
D27090 N27090 0 diode
R27091 N27090 N27091 10
D27091 N27091 0 diode
R27092 N27091 N27092 10
D27092 N27092 0 diode
R27093 N27092 N27093 10
D27093 N27093 0 diode
R27094 N27093 N27094 10
D27094 N27094 0 diode
R27095 N27094 N27095 10
D27095 N27095 0 diode
R27096 N27095 N27096 10
D27096 N27096 0 diode
R27097 N27096 N27097 10
D27097 N27097 0 diode
R27098 N27097 N27098 10
D27098 N27098 0 diode
R27099 N27098 N27099 10
D27099 N27099 0 diode
R27100 N27099 N27100 10
D27100 N27100 0 diode
R27101 N27100 N27101 10
D27101 N27101 0 diode
R27102 N27101 N27102 10
D27102 N27102 0 diode
R27103 N27102 N27103 10
D27103 N27103 0 diode
R27104 N27103 N27104 10
D27104 N27104 0 diode
R27105 N27104 N27105 10
D27105 N27105 0 diode
R27106 N27105 N27106 10
D27106 N27106 0 diode
R27107 N27106 N27107 10
D27107 N27107 0 diode
R27108 N27107 N27108 10
D27108 N27108 0 diode
R27109 N27108 N27109 10
D27109 N27109 0 diode
R27110 N27109 N27110 10
D27110 N27110 0 diode
R27111 N27110 N27111 10
D27111 N27111 0 diode
R27112 N27111 N27112 10
D27112 N27112 0 diode
R27113 N27112 N27113 10
D27113 N27113 0 diode
R27114 N27113 N27114 10
D27114 N27114 0 diode
R27115 N27114 N27115 10
D27115 N27115 0 diode
R27116 N27115 N27116 10
D27116 N27116 0 diode
R27117 N27116 N27117 10
D27117 N27117 0 diode
R27118 N27117 N27118 10
D27118 N27118 0 diode
R27119 N27118 N27119 10
D27119 N27119 0 diode
R27120 N27119 N27120 10
D27120 N27120 0 diode
R27121 N27120 N27121 10
D27121 N27121 0 diode
R27122 N27121 N27122 10
D27122 N27122 0 diode
R27123 N27122 N27123 10
D27123 N27123 0 diode
R27124 N27123 N27124 10
D27124 N27124 0 diode
R27125 N27124 N27125 10
D27125 N27125 0 diode
R27126 N27125 N27126 10
D27126 N27126 0 diode
R27127 N27126 N27127 10
D27127 N27127 0 diode
R27128 N27127 N27128 10
D27128 N27128 0 diode
R27129 N27128 N27129 10
D27129 N27129 0 diode
R27130 N27129 N27130 10
D27130 N27130 0 diode
R27131 N27130 N27131 10
D27131 N27131 0 diode
R27132 N27131 N27132 10
D27132 N27132 0 diode
R27133 N27132 N27133 10
D27133 N27133 0 diode
R27134 N27133 N27134 10
D27134 N27134 0 diode
R27135 N27134 N27135 10
D27135 N27135 0 diode
R27136 N27135 N27136 10
D27136 N27136 0 diode
R27137 N27136 N27137 10
D27137 N27137 0 diode
R27138 N27137 N27138 10
D27138 N27138 0 diode
R27139 N27138 N27139 10
D27139 N27139 0 diode
R27140 N27139 N27140 10
D27140 N27140 0 diode
R27141 N27140 N27141 10
D27141 N27141 0 diode
R27142 N27141 N27142 10
D27142 N27142 0 diode
R27143 N27142 N27143 10
D27143 N27143 0 diode
R27144 N27143 N27144 10
D27144 N27144 0 diode
R27145 N27144 N27145 10
D27145 N27145 0 diode
R27146 N27145 N27146 10
D27146 N27146 0 diode
R27147 N27146 N27147 10
D27147 N27147 0 diode
R27148 N27147 N27148 10
D27148 N27148 0 diode
R27149 N27148 N27149 10
D27149 N27149 0 diode
R27150 N27149 N27150 10
D27150 N27150 0 diode
R27151 N27150 N27151 10
D27151 N27151 0 diode
R27152 N27151 N27152 10
D27152 N27152 0 diode
R27153 N27152 N27153 10
D27153 N27153 0 diode
R27154 N27153 N27154 10
D27154 N27154 0 diode
R27155 N27154 N27155 10
D27155 N27155 0 diode
R27156 N27155 N27156 10
D27156 N27156 0 diode
R27157 N27156 N27157 10
D27157 N27157 0 diode
R27158 N27157 N27158 10
D27158 N27158 0 diode
R27159 N27158 N27159 10
D27159 N27159 0 diode
R27160 N27159 N27160 10
D27160 N27160 0 diode
R27161 N27160 N27161 10
D27161 N27161 0 diode
R27162 N27161 N27162 10
D27162 N27162 0 diode
R27163 N27162 N27163 10
D27163 N27163 0 diode
R27164 N27163 N27164 10
D27164 N27164 0 diode
R27165 N27164 N27165 10
D27165 N27165 0 diode
R27166 N27165 N27166 10
D27166 N27166 0 diode
R27167 N27166 N27167 10
D27167 N27167 0 diode
R27168 N27167 N27168 10
D27168 N27168 0 diode
R27169 N27168 N27169 10
D27169 N27169 0 diode
R27170 N27169 N27170 10
D27170 N27170 0 diode
R27171 N27170 N27171 10
D27171 N27171 0 diode
R27172 N27171 N27172 10
D27172 N27172 0 diode
R27173 N27172 N27173 10
D27173 N27173 0 diode
R27174 N27173 N27174 10
D27174 N27174 0 diode
R27175 N27174 N27175 10
D27175 N27175 0 diode
R27176 N27175 N27176 10
D27176 N27176 0 diode
R27177 N27176 N27177 10
D27177 N27177 0 diode
R27178 N27177 N27178 10
D27178 N27178 0 diode
R27179 N27178 N27179 10
D27179 N27179 0 diode
R27180 N27179 N27180 10
D27180 N27180 0 diode
R27181 N27180 N27181 10
D27181 N27181 0 diode
R27182 N27181 N27182 10
D27182 N27182 0 diode
R27183 N27182 N27183 10
D27183 N27183 0 diode
R27184 N27183 N27184 10
D27184 N27184 0 diode
R27185 N27184 N27185 10
D27185 N27185 0 diode
R27186 N27185 N27186 10
D27186 N27186 0 diode
R27187 N27186 N27187 10
D27187 N27187 0 diode
R27188 N27187 N27188 10
D27188 N27188 0 diode
R27189 N27188 N27189 10
D27189 N27189 0 diode
R27190 N27189 N27190 10
D27190 N27190 0 diode
R27191 N27190 N27191 10
D27191 N27191 0 diode
R27192 N27191 N27192 10
D27192 N27192 0 diode
R27193 N27192 N27193 10
D27193 N27193 0 diode
R27194 N27193 N27194 10
D27194 N27194 0 diode
R27195 N27194 N27195 10
D27195 N27195 0 diode
R27196 N27195 N27196 10
D27196 N27196 0 diode
R27197 N27196 N27197 10
D27197 N27197 0 diode
R27198 N27197 N27198 10
D27198 N27198 0 diode
R27199 N27198 N27199 10
D27199 N27199 0 diode
R27200 N27199 N27200 10
D27200 N27200 0 diode
R27201 N27200 N27201 10
D27201 N27201 0 diode
R27202 N27201 N27202 10
D27202 N27202 0 diode
R27203 N27202 N27203 10
D27203 N27203 0 diode
R27204 N27203 N27204 10
D27204 N27204 0 diode
R27205 N27204 N27205 10
D27205 N27205 0 diode
R27206 N27205 N27206 10
D27206 N27206 0 diode
R27207 N27206 N27207 10
D27207 N27207 0 diode
R27208 N27207 N27208 10
D27208 N27208 0 diode
R27209 N27208 N27209 10
D27209 N27209 0 diode
R27210 N27209 N27210 10
D27210 N27210 0 diode
R27211 N27210 N27211 10
D27211 N27211 0 diode
R27212 N27211 N27212 10
D27212 N27212 0 diode
R27213 N27212 N27213 10
D27213 N27213 0 diode
R27214 N27213 N27214 10
D27214 N27214 0 diode
R27215 N27214 N27215 10
D27215 N27215 0 diode
R27216 N27215 N27216 10
D27216 N27216 0 diode
R27217 N27216 N27217 10
D27217 N27217 0 diode
R27218 N27217 N27218 10
D27218 N27218 0 diode
R27219 N27218 N27219 10
D27219 N27219 0 diode
R27220 N27219 N27220 10
D27220 N27220 0 diode
R27221 N27220 N27221 10
D27221 N27221 0 diode
R27222 N27221 N27222 10
D27222 N27222 0 diode
R27223 N27222 N27223 10
D27223 N27223 0 diode
R27224 N27223 N27224 10
D27224 N27224 0 diode
R27225 N27224 N27225 10
D27225 N27225 0 diode
R27226 N27225 N27226 10
D27226 N27226 0 diode
R27227 N27226 N27227 10
D27227 N27227 0 diode
R27228 N27227 N27228 10
D27228 N27228 0 diode
R27229 N27228 N27229 10
D27229 N27229 0 diode
R27230 N27229 N27230 10
D27230 N27230 0 diode
R27231 N27230 N27231 10
D27231 N27231 0 diode
R27232 N27231 N27232 10
D27232 N27232 0 diode
R27233 N27232 N27233 10
D27233 N27233 0 diode
R27234 N27233 N27234 10
D27234 N27234 0 diode
R27235 N27234 N27235 10
D27235 N27235 0 diode
R27236 N27235 N27236 10
D27236 N27236 0 diode
R27237 N27236 N27237 10
D27237 N27237 0 diode
R27238 N27237 N27238 10
D27238 N27238 0 diode
R27239 N27238 N27239 10
D27239 N27239 0 diode
R27240 N27239 N27240 10
D27240 N27240 0 diode
R27241 N27240 N27241 10
D27241 N27241 0 diode
R27242 N27241 N27242 10
D27242 N27242 0 diode
R27243 N27242 N27243 10
D27243 N27243 0 diode
R27244 N27243 N27244 10
D27244 N27244 0 diode
R27245 N27244 N27245 10
D27245 N27245 0 diode
R27246 N27245 N27246 10
D27246 N27246 0 diode
R27247 N27246 N27247 10
D27247 N27247 0 diode
R27248 N27247 N27248 10
D27248 N27248 0 diode
R27249 N27248 N27249 10
D27249 N27249 0 diode
R27250 N27249 N27250 10
D27250 N27250 0 diode
R27251 N27250 N27251 10
D27251 N27251 0 diode
R27252 N27251 N27252 10
D27252 N27252 0 diode
R27253 N27252 N27253 10
D27253 N27253 0 diode
R27254 N27253 N27254 10
D27254 N27254 0 diode
R27255 N27254 N27255 10
D27255 N27255 0 diode
R27256 N27255 N27256 10
D27256 N27256 0 diode
R27257 N27256 N27257 10
D27257 N27257 0 diode
R27258 N27257 N27258 10
D27258 N27258 0 diode
R27259 N27258 N27259 10
D27259 N27259 0 diode
R27260 N27259 N27260 10
D27260 N27260 0 diode
R27261 N27260 N27261 10
D27261 N27261 0 diode
R27262 N27261 N27262 10
D27262 N27262 0 diode
R27263 N27262 N27263 10
D27263 N27263 0 diode
R27264 N27263 N27264 10
D27264 N27264 0 diode
R27265 N27264 N27265 10
D27265 N27265 0 diode
R27266 N27265 N27266 10
D27266 N27266 0 diode
R27267 N27266 N27267 10
D27267 N27267 0 diode
R27268 N27267 N27268 10
D27268 N27268 0 diode
R27269 N27268 N27269 10
D27269 N27269 0 diode
R27270 N27269 N27270 10
D27270 N27270 0 diode
R27271 N27270 N27271 10
D27271 N27271 0 diode
R27272 N27271 N27272 10
D27272 N27272 0 diode
R27273 N27272 N27273 10
D27273 N27273 0 diode
R27274 N27273 N27274 10
D27274 N27274 0 diode
R27275 N27274 N27275 10
D27275 N27275 0 diode
R27276 N27275 N27276 10
D27276 N27276 0 diode
R27277 N27276 N27277 10
D27277 N27277 0 diode
R27278 N27277 N27278 10
D27278 N27278 0 diode
R27279 N27278 N27279 10
D27279 N27279 0 diode
R27280 N27279 N27280 10
D27280 N27280 0 diode
R27281 N27280 N27281 10
D27281 N27281 0 diode
R27282 N27281 N27282 10
D27282 N27282 0 diode
R27283 N27282 N27283 10
D27283 N27283 0 diode
R27284 N27283 N27284 10
D27284 N27284 0 diode
R27285 N27284 N27285 10
D27285 N27285 0 diode
R27286 N27285 N27286 10
D27286 N27286 0 diode
R27287 N27286 N27287 10
D27287 N27287 0 diode
R27288 N27287 N27288 10
D27288 N27288 0 diode
R27289 N27288 N27289 10
D27289 N27289 0 diode
R27290 N27289 N27290 10
D27290 N27290 0 diode
R27291 N27290 N27291 10
D27291 N27291 0 diode
R27292 N27291 N27292 10
D27292 N27292 0 diode
R27293 N27292 N27293 10
D27293 N27293 0 diode
R27294 N27293 N27294 10
D27294 N27294 0 diode
R27295 N27294 N27295 10
D27295 N27295 0 diode
R27296 N27295 N27296 10
D27296 N27296 0 diode
R27297 N27296 N27297 10
D27297 N27297 0 diode
R27298 N27297 N27298 10
D27298 N27298 0 diode
R27299 N27298 N27299 10
D27299 N27299 0 diode
R27300 N27299 N27300 10
D27300 N27300 0 diode
R27301 N27300 N27301 10
D27301 N27301 0 diode
R27302 N27301 N27302 10
D27302 N27302 0 diode
R27303 N27302 N27303 10
D27303 N27303 0 diode
R27304 N27303 N27304 10
D27304 N27304 0 diode
R27305 N27304 N27305 10
D27305 N27305 0 diode
R27306 N27305 N27306 10
D27306 N27306 0 diode
R27307 N27306 N27307 10
D27307 N27307 0 diode
R27308 N27307 N27308 10
D27308 N27308 0 diode
R27309 N27308 N27309 10
D27309 N27309 0 diode
R27310 N27309 N27310 10
D27310 N27310 0 diode
R27311 N27310 N27311 10
D27311 N27311 0 diode
R27312 N27311 N27312 10
D27312 N27312 0 diode
R27313 N27312 N27313 10
D27313 N27313 0 diode
R27314 N27313 N27314 10
D27314 N27314 0 diode
R27315 N27314 N27315 10
D27315 N27315 0 diode
R27316 N27315 N27316 10
D27316 N27316 0 diode
R27317 N27316 N27317 10
D27317 N27317 0 diode
R27318 N27317 N27318 10
D27318 N27318 0 diode
R27319 N27318 N27319 10
D27319 N27319 0 diode
R27320 N27319 N27320 10
D27320 N27320 0 diode
R27321 N27320 N27321 10
D27321 N27321 0 diode
R27322 N27321 N27322 10
D27322 N27322 0 diode
R27323 N27322 N27323 10
D27323 N27323 0 diode
R27324 N27323 N27324 10
D27324 N27324 0 diode
R27325 N27324 N27325 10
D27325 N27325 0 diode
R27326 N27325 N27326 10
D27326 N27326 0 diode
R27327 N27326 N27327 10
D27327 N27327 0 diode
R27328 N27327 N27328 10
D27328 N27328 0 diode
R27329 N27328 N27329 10
D27329 N27329 0 diode
R27330 N27329 N27330 10
D27330 N27330 0 diode
R27331 N27330 N27331 10
D27331 N27331 0 diode
R27332 N27331 N27332 10
D27332 N27332 0 diode
R27333 N27332 N27333 10
D27333 N27333 0 diode
R27334 N27333 N27334 10
D27334 N27334 0 diode
R27335 N27334 N27335 10
D27335 N27335 0 diode
R27336 N27335 N27336 10
D27336 N27336 0 diode
R27337 N27336 N27337 10
D27337 N27337 0 diode
R27338 N27337 N27338 10
D27338 N27338 0 diode
R27339 N27338 N27339 10
D27339 N27339 0 diode
R27340 N27339 N27340 10
D27340 N27340 0 diode
R27341 N27340 N27341 10
D27341 N27341 0 diode
R27342 N27341 N27342 10
D27342 N27342 0 diode
R27343 N27342 N27343 10
D27343 N27343 0 diode
R27344 N27343 N27344 10
D27344 N27344 0 diode
R27345 N27344 N27345 10
D27345 N27345 0 diode
R27346 N27345 N27346 10
D27346 N27346 0 diode
R27347 N27346 N27347 10
D27347 N27347 0 diode
R27348 N27347 N27348 10
D27348 N27348 0 diode
R27349 N27348 N27349 10
D27349 N27349 0 diode
R27350 N27349 N27350 10
D27350 N27350 0 diode
R27351 N27350 N27351 10
D27351 N27351 0 diode
R27352 N27351 N27352 10
D27352 N27352 0 diode
R27353 N27352 N27353 10
D27353 N27353 0 diode
R27354 N27353 N27354 10
D27354 N27354 0 diode
R27355 N27354 N27355 10
D27355 N27355 0 diode
R27356 N27355 N27356 10
D27356 N27356 0 diode
R27357 N27356 N27357 10
D27357 N27357 0 diode
R27358 N27357 N27358 10
D27358 N27358 0 diode
R27359 N27358 N27359 10
D27359 N27359 0 diode
R27360 N27359 N27360 10
D27360 N27360 0 diode
R27361 N27360 N27361 10
D27361 N27361 0 diode
R27362 N27361 N27362 10
D27362 N27362 0 diode
R27363 N27362 N27363 10
D27363 N27363 0 diode
R27364 N27363 N27364 10
D27364 N27364 0 diode
R27365 N27364 N27365 10
D27365 N27365 0 diode
R27366 N27365 N27366 10
D27366 N27366 0 diode
R27367 N27366 N27367 10
D27367 N27367 0 diode
R27368 N27367 N27368 10
D27368 N27368 0 diode
R27369 N27368 N27369 10
D27369 N27369 0 diode
R27370 N27369 N27370 10
D27370 N27370 0 diode
R27371 N27370 N27371 10
D27371 N27371 0 diode
R27372 N27371 N27372 10
D27372 N27372 0 diode
R27373 N27372 N27373 10
D27373 N27373 0 diode
R27374 N27373 N27374 10
D27374 N27374 0 diode
R27375 N27374 N27375 10
D27375 N27375 0 diode
R27376 N27375 N27376 10
D27376 N27376 0 diode
R27377 N27376 N27377 10
D27377 N27377 0 diode
R27378 N27377 N27378 10
D27378 N27378 0 diode
R27379 N27378 N27379 10
D27379 N27379 0 diode
R27380 N27379 N27380 10
D27380 N27380 0 diode
R27381 N27380 N27381 10
D27381 N27381 0 diode
R27382 N27381 N27382 10
D27382 N27382 0 diode
R27383 N27382 N27383 10
D27383 N27383 0 diode
R27384 N27383 N27384 10
D27384 N27384 0 diode
R27385 N27384 N27385 10
D27385 N27385 0 diode
R27386 N27385 N27386 10
D27386 N27386 0 diode
R27387 N27386 N27387 10
D27387 N27387 0 diode
R27388 N27387 N27388 10
D27388 N27388 0 diode
R27389 N27388 N27389 10
D27389 N27389 0 diode
R27390 N27389 N27390 10
D27390 N27390 0 diode
R27391 N27390 N27391 10
D27391 N27391 0 diode
R27392 N27391 N27392 10
D27392 N27392 0 diode
R27393 N27392 N27393 10
D27393 N27393 0 diode
R27394 N27393 N27394 10
D27394 N27394 0 diode
R27395 N27394 N27395 10
D27395 N27395 0 diode
R27396 N27395 N27396 10
D27396 N27396 0 diode
R27397 N27396 N27397 10
D27397 N27397 0 diode
R27398 N27397 N27398 10
D27398 N27398 0 diode
R27399 N27398 N27399 10
D27399 N27399 0 diode
R27400 N27399 N27400 10
D27400 N27400 0 diode
R27401 N27400 N27401 10
D27401 N27401 0 diode
R27402 N27401 N27402 10
D27402 N27402 0 diode
R27403 N27402 N27403 10
D27403 N27403 0 diode
R27404 N27403 N27404 10
D27404 N27404 0 diode
R27405 N27404 N27405 10
D27405 N27405 0 diode
R27406 N27405 N27406 10
D27406 N27406 0 diode
R27407 N27406 N27407 10
D27407 N27407 0 diode
R27408 N27407 N27408 10
D27408 N27408 0 diode
R27409 N27408 N27409 10
D27409 N27409 0 diode
R27410 N27409 N27410 10
D27410 N27410 0 diode
R27411 N27410 N27411 10
D27411 N27411 0 diode
R27412 N27411 N27412 10
D27412 N27412 0 diode
R27413 N27412 N27413 10
D27413 N27413 0 diode
R27414 N27413 N27414 10
D27414 N27414 0 diode
R27415 N27414 N27415 10
D27415 N27415 0 diode
R27416 N27415 N27416 10
D27416 N27416 0 diode
R27417 N27416 N27417 10
D27417 N27417 0 diode
R27418 N27417 N27418 10
D27418 N27418 0 diode
R27419 N27418 N27419 10
D27419 N27419 0 diode
R27420 N27419 N27420 10
D27420 N27420 0 diode
R27421 N27420 N27421 10
D27421 N27421 0 diode
R27422 N27421 N27422 10
D27422 N27422 0 diode
R27423 N27422 N27423 10
D27423 N27423 0 diode
R27424 N27423 N27424 10
D27424 N27424 0 diode
R27425 N27424 N27425 10
D27425 N27425 0 diode
R27426 N27425 N27426 10
D27426 N27426 0 diode
R27427 N27426 N27427 10
D27427 N27427 0 diode
R27428 N27427 N27428 10
D27428 N27428 0 diode
R27429 N27428 N27429 10
D27429 N27429 0 diode
R27430 N27429 N27430 10
D27430 N27430 0 diode
R27431 N27430 N27431 10
D27431 N27431 0 diode
R27432 N27431 N27432 10
D27432 N27432 0 diode
R27433 N27432 N27433 10
D27433 N27433 0 diode
R27434 N27433 N27434 10
D27434 N27434 0 diode
R27435 N27434 N27435 10
D27435 N27435 0 diode
R27436 N27435 N27436 10
D27436 N27436 0 diode
R27437 N27436 N27437 10
D27437 N27437 0 diode
R27438 N27437 N27438 10
D27438 N27438 0 diode
R27439 N27438 N27439 10
D27439 N27439 0 diode
R27440 N27439 N27440 10
D27440 N27440 0 diode
R27441 N27440 N27441 10
D27441 N27441 0 diode
R27442 N27441 N27442 10
D27442 N27442 0 diode
R27443 N27442 N27443 10
D27443 N27443 0 diode
R27444 N27443 N27444 10
D27444 N27444 0 diode
R27445 N27444 N27445 10
D27445 N27445 0 diode
R27446 N27445 N27446 10
D27446 N27446 0 diode
R27447 N27446 N27447 10
D27447 N27447 0 diode
R27448 N27447 N27448 10
D27448 N27448 0 diode
R27449 N27448 N27449 10
D27449 N27449 0 diode
R27450 N27449 N27450 10
D27450 N27450 0 diode
R27451 N27450 N27451 10
D27451 N27451 0 diode
R27452 N27451 N27452 10
D27452 N27452 0 diode
R27453 N27452 N27453 10
D27453 N27453 0 diode
R27454 N27453 N27454 10
D27454 N27454 0 diode
R27455 N27454 N27455 10
D27455 N27455 0 diode
R27456 N27455 N27456 10
D27456 N27456 0 diode
R27457 N27456 N27457 10
D27457 N27457 0 diode
R27458 N27457 N27458 10
D27458 N27458 0 diode
R27459 N27458 N27459 10
D27459 N27459 0 diode
R27460 N27459 N27460 10
D27460 N27460 0 diode
R27461 N27460 N27461 10
D27461 N27461 0 diode
R27462 N27461 N27462 10
D27462 N27462 0 diode
R27463 N27462 N27463 10
D27463 N27463 0 diode
R27464 N27463 N27464 10
D27464 N27464 0 diode
R27465 N27464 N27465 10
D27465 N27465 0 diode
R27466 N27465 N27466 10
D27466 N27466 0 diode
R27467 N27466 N27467 10
D27467 N27467 0 diode
R27468 N27467 N27468 10
D27468 N27468 0 diode
R27469 N27468 N27469 10
D27469 N27469 0 diode
R27470 N27469 N27470 10
D27470 N27470 0 diode
R27471 N27470 N27471 10
D27471 N27471 0 diode
R27472 N27471 N27472 10
D27472 N27472 0 diode
R27473 N27472 N27473 10
D27473 N27473 0 diode
R27474 N27473 N27474 10
D27474 N27474 0 diode
R27475 N27474 N27475 10
D27475 N27475 0 diode
R27476 N27475 N27476 10
D27476 N27476 0 diode
R27477 N27476 N27477 10
D27477 N27477 0 diode
R27478 N27477 N27478 10
D27478 N27478 0 diode
R27479 N27478 N27479 10
D27479 N27479 0 diode
R27480 N27479 N27480 10
D27480 N27480 0 diode
R27481 N27480 N27481 10
D27481 N27481 0 diode
R27482 N27481 N27482 10
D27482 N27482 0 diode
R27483 N27482 N27483 10
D27483 N27483 0 diode
R27484 N27483 N27484 10
D27484 N27484 0 diode
R27485 N27484 N27485 10
D27485 N27485 0 diode
R27486 N27485 N27486 10
D27486 N27486 0 diode
R27487 N27486 N27487 10
D27487 N27487 0 diode
R27488 N27487 N27488 10
D27488 N27488 0 diode
R27489 N27488 N27489 10
D27489 N27489 0 diode
R27490 N27489 N27490 10
D27490 N27490 0 diode
R27491 N27490 N27491 10
D27491 N27491 0 diode
R27492 N27491 N27492 10
D27492 N27492 0 diode
R27493 N27492 N27493 10
D27493 N27493 0 diode
R27494 N27493 N27494 10
D27494 N27494 0 diode
R27495 N27494 N27495 10
D27495 N27495 0 diode
R27496 N27495 N27496 10
D27496 N27496 0 diode
R27497 N27496 N27497 10
D27497 N27497 0 diode
R27498 N27497 N27498 10
D27498 N27498 0 diode
R27499 N27498 N27499 10
D27499 N27499 0 diode
R27500 N27499 N27500 10
D27500 N27500 0 diode
R27501 N27500 N27501 10
D27501 N27501 0 diode
R27502 N27501 N27502 10
D27502 N27502 0 diode
R27503 N27502 N27503 10
D27503 N27503 0 diode
R27504 N27503 N27504 10
D27504 N27504 0 diode
R27505 N27504 N27505 10
D27505 N27505 0 diode
R27506 N27505 N27506 10
D27506 N27506 0 diode
R27507 N27506 N27507 10
D27507 N27507 0 diode
R27508 N27507 N27508 10
D27508 N27508 0 diode
R27509 N27508 N27509 10
D27509 N27509 0 diode
R27510 N27509 N27510 10
D27510 N27510 0 diode
R27511 N27510 N27511 10
D27511 N27511 0 diode
R27512 N27511 N27512 10
D27512 N27512 0 diode
R27513 N27512 N27513 10
D27513 N27513 0 diode
R27514 N27513 N27514 10
D27514 N27514 0 diode
R27515 N27514 N27515 10
D27515 N27515 0 diode
R27516 N27515 N27516 10
D27516 N27516 0 diode
R27517 N27516 N27517 10
D27517 N27517 0 diode
R27518 N27517 N27518 10
D27518 N27518 0 diode
R27519 N27518 N27519 10
D27519 N27519 0 diode
R27520 N27519 N27520 10
D27520 N27520 0 diode
R27521 N27520 N27521 10
D27521 N27521 0 diode
R27522 N27521 N27522 10
D27522 N27522 0 diode
R27523 N27522 N27523 10
D27523 N27523 0 diode
R27524 N27523 N27524 10
D27524 N27524 0 diode
R27525 N27524 N27525 10
D27525 N27525 0 diode
R27526 N27525 N27526 10
D27526 N27526 0 diode
R27527 N27526 N27527 10
D27527 N27527 0 diode
R27528 N27527 N27528 10
D27528 N27528 0 diode
R27529 N27528 N27529 10
D27529 N27529 0 diode
R27530 N27529 N27530 10
D27530 N27530 0 diode
R27531 N27530 N27531 10
D27531 N27531 0 diode
R27532 N27531 N27532 10
D27532 N27532 0 diode
R27533 N27532 N27533 10
D27533 N27533 0 diode
R27534 N27533 N27534 10
D27534 N27534 0 diode
R27535 N27534 N27535 10
D27535 N27535 0 diode
R27536 N27535 N27536 10
D27536 N27536 0 diode
R27537 N27536 N27537 10
D27537 N27537 0 diode
R27538 N27537 N27538 10
D27538 N27538 0 diode
R27539 N27538 N27539 10
D27539 N27539 0 diode
R27540 N27539 N27540 10
D27540 N27540 0 diode
R27541 N27540 N27541 10
D27541 N27541 0 diode
R27542 N27541 N27542 10
D27542 N27542 0 diode
R27543 N27542 N27543 10
D27543 N27543 0 diode
R27544 N27543 N27544 10
D27544 N27544 0 diode
R27545 N27544 N27545 10
D27545 N27545 0 diode
R27546 N27545 N27546 10
D27546 N27546 0 diode
R27547 N27546 N27547 10
D27547 N27547 0 diode
R27548 N27547 N27548 10
D27548 N27548 0 diode
R27549 N27548 N27549 10
D27549 N27549 0 diode
R27550 N27549 N27550 10
D27550 N27550 0 diode
R27551 N27550 N27551 10
D27551 N27551 0 diode
R27552 N27551 N27552 10
D27552 N27552 0 diode
R27553 N27552 N27553 10
D27553 N27553 0 diode
R27554 N27553 N27554 10
D27554 N27554 0 diode
R27555 N27554 N27555 10
D27555 N27555 0 diode
R27556 N27555 N27556 10
D27556 N27556 0 diode
R27557 N27556 N27557 10
D27557 N27557 0 diode
R27558 N27557 N27558 10
D27558 N27558 0 diode
R27559 N27558 N27559 10
D27559 N27559 0 diode
R27560 N27559 N27560 10
D27560 N27560 0 diode
R27561 N27560 N27561 10
D27561 N27561 0 diode
R27562 N27561 N27562 10
D27562 N27562 0 diode
R27563 N27562 N27563 10
D27563 N27563 0 diode
R27564 N27563 N27564 10
D27564 N27564 0 diode
R27565 N27564 N27565 10
D27565 N27565 0 diode
R27566 N27565 N27566 10
D27566 N27566 0 diode
R27567 N27566 N27567 10
D27567 N27567 0 diode
R27568 N27567 N27568 10
D27568 N27568 0 diode
R27569 N27568 N27569 10
D27569 N27569 0 diode
R27570 N27569 N27570 10
D27570 N27570 0 diode
R27571 N27570 N27571 10
D27571 N27571 0 diode
R27572 N27571 N27572 10
D27572 N27572 0 diode
R27573 N27572 N27573 10
D27573 N27573 0 diode
R27574 N27573 N27574 10
D27574 N27574 0 diode
R27575 N27574 N27575 10
D27575 N27575 0 diode
R27576 N27575 N27576 10
D27576 N27576 0 diode
R27577 N27576 N27577 10
D27577 N27577 0 diode
R27578 N27577 N27578 10
D27578 N27578 0 diode
R27579 N27578 N27579 10
D27579 N27579 0 diode
R27580 N27579 N27580 10
D27580 N27580 0 diode
R27581 N27580 N27581 10
D27581 N27581 0 diode
R27582 N27581 N27582 10
D27582 N27582 0 diode
R27583 N27582 N27583 10
D27583 N27583 0 diode
R27584 N27583 N27584 10
D27584 N27584 0 diode
R27585 N27584 N27585 10
D27585 N27585 0 diode
R27586 N27585 N27586 10
D27586 N27586 0 diode
R27587 N27586 N27587 10
D27587 N27587 0 diode
R27588 N27587 N27588 10
D27588 N27588 0 diode
R27589 N27588 N27589 10
D27589 N27589 0 diode
R27590 N27589 N27590 10
D27590 N27590 0 diode
R27591 N27590 N27591 10
D27591 N27591 0 diode
R27592 N27591 N27592 10
D27592 N27592 0 diode
R27593 N27592 N27593 10
D27593 N27593 0 diode
R27594 N27593 N27594 10
D27594 N27594 0 diode
R27595 N27594 N27595 10
D27595 N27595 0 diode
R27596 N27595 N27596 10
D27596 N27596 0 diode
R27597 N27596 N27597 10
D27597 N27597 0 diode
R27598 N27597 N27598 10
D27598 N27598 0 diode
R27599 N27598 N27599 10
D27599 N27599 0 diode
R27600 N27599 N27600 10
D27600 N27600 0 diode
R27601 N27600 N27601 10
D27601 N27601 0 diode
R27602 N27601 N27602 10
D27602 N27602 0 diode
R27603 N27602 N27603 10
D27603 N27603 0 diode
R27604 N27603 N27604 10
D27604 N27604 0 diode
R27605 N27604 N27605 10
D27605 N27605 0 diode
R27606 N27605 N27606 10
D27606 N27606 0 diode
R27607 N27606 N27607 10
D27607 N27607 0 diode
R27608 N27607 N27608 10
D27608 N27608 0 diode
R27609 N27608 N27609 10
D27609 N27609 0 diode
R27610 N27609 N27610 10
D27610 N27610 0 diode
R27611 N27610 N27611 10
D27611 N27611 0 diode
R27612 N27611 N27612 10
D27612 N27612 0 diode
R27613 N27612 N27613 10
D27613 N27613 0 diode
R27614 N27613 N27614 10
D27614 N27614 0 diode
R27615 N27614 N27615 10
D27615 N27615 0 diode
R27616 N27615 N27616 10
D27616 N27616 0 diode
R27617 N27616 N27617 10
D27617 N27617 0 diode
R27618 N27617 N27618 10
D27618 N27618 0 diode
R27619 N27618 N27619 10
D27619 N27619 0 diode
R27620 N27619 N27620 10
D27620 N27620 0 diode
R27621 N27620 N27621 10
D27621 N27621 0 diode
R27622 N27621 N27622 10
D27622 N27622 0 diode
R27623 N27622 N27623 10
D27623 N27623 0 diode
R27624 N27623 N27624 10
D27624 N27624 0 diode
R27625 N27624 N27625 10
D27625 N27625 0 diode
R27626 N27625 N27626 10
D27626 N27626 0 diode
R27627 N27626 N27627 10
D27627 N27627 0 diode
R27628 N27627 N27628 10
D27628 N27628 0 diode
R27629 N27628 N27629 10
D27629 N27629 0 diode
R27630 N27629 N27630 10
D27630 N27630 0 diode
R27631 N27630 N27631 10
D27631 N27631 0 diode
R27632 N27631 N27632 10
D27632 N27632 0 diode
R27633 N27632 N27633 10
D27633 N27633 0 diode
R27634 N27633 N27634 10
D27634 N27634 0 diode
R27635 N27634 N27635 10
D27635 N27635 0 diode
R27636 N27635 N27636 10
D27636 N27636 0 diode
R27637 N27636 N27637 10
D27637 N27637 0 diode
R27638 N27637 N27638 10
D27638 N27638 0 diode
R27639 N27638 N27639 10
D27639 N27639 0 diode
R27640 N27639 N27640 10
D27640 N27640 0 diode
R27641 N27640 N27641 10
D27641 N27641 0 diode
R27642 N27641 N27642 10
D27642 N27642 0 diode
R27643 N27642 N27643 10
D27643 N27643 0 diode
R27644 N27643 N27644 10
D27644 N27644 0 diode
R27645 N27644 N27645 10
D27645 N27645 0 diode
R27646 N27645 N27646 10
D27646 N27646 0 diode
R27647 N27646 N27647 10
D27647 N27647 0 diode
R27648 N27647 N27648 10
D27648 N27648 0 diode
R27649 N27648 N27649 10
D27649 N27649 0 diode
R27650 N27649 N27650 10
D27650 N27650 0 diode
R27651 N27650 N27651 10
D27651 N27651 0 diode
R27652 N27651 N27652 10
D27652 N27652 0 diode
R27653 N27652 N27653 10
D27653 N27653 0 diode
R27654 N27653 N27654 10
D27654 N27654 0 diode
R27655 N27654 N27655 10
D27655 N27655 0 diode
R27656 N27655 N27656 10
D27656 N27656 0 diode
R27657 N27656 N27657 10
D27657 N27657 0 diode
R27658 N27657 N27658 10
D27658 N27658 0 diode
R27659 N27658 N27659 10
D27659 N27659 0 diode
R27660 N27659 N27660 10
D27660 N27660 0 diode
R27661 N27660 N27661 10
D27661 N27661 0 diode
R27662 N27661 N27662 10
D27662 N27662 0 diode
R27663 N27662 N27663 10
D27663 N27663 0 diode
R27664 N27663 N27664 10
D27664 N27664 0 diode
R27665 N27664 N27665 10
D27665 N27665 0 diode
R27666 N27665 N27666 10
D27666 N27666 0 diode
R27667 N27666 N27667 10
D27667 N27667 0 diode
R27668 N27667 N27668 10
D27668 N27668 0 diode
R27669 N27668 N27669 10
D27669 N27669 0 diode
R27670 N27669 N27670 10
D27670 N27670 0 diode
R27671 N27670 N27671 10
D27671 N27671 0 diode
R27672 N27671 N27672 10
D27672 N27672 0 diode
R27673 N27672 N27673 10
D27673 N27673 0 diode
R27674 N27673 N27674 10
D27674 N27674 0 diode
R27675 N27674 N27675 10
D27675 N27675 0 diode
R27676 N27675 N27676 10
D27676 N27676 0 diode
R27677 N27676 N27677 10
D27677 N27677 0 diode
R27678 N27677 N27678 10
D27678 N27678 0 diode
R27679 N27678 N27679 10
D27679 N27679 0 diode
R27680 N27679 N27680 10
D27680 N27680 0 diode
R27681 N27680 N27681 10
D27681 N27681 0 diode
R27682 N27681 N27682 10
D27682 N27682 0 diode
R27683 N27682 N27683 10
D27683 N27683 0 diode
R27684 N27683 N27684 10
D27684 N27684 0 diode
R27685 N27684 N27685 10
D27685 N27685 0 diode
R27686 N27685 N27686 10
D27686 N27686 0 diode
R27687 N27686 N27687 10
D27687 N27687 0 diode
R27688 N27687 N27688 10
D27688 N27688 0 diode
R27689 N27688 N27689 10
D27689 N27689 0 diode
R27690 N27689 N27690 10
D27690 N27690 0 diode
R27691 N27690 N27691 10
D27691 N27691 0 diode
R27692 N27691 N27692 10
D27692 N27692 0 diode
R27693 N27692 N27693 10
D27693 N27693 0 diode
R27694 N27693 N27694 10
D27694 N27694 0 diode
R27695 N27694 N27695 10
D27695 N27695 0 diode
R27696 N27695 N27696 10
D27696 N27696 0 diode
R27697 N27696 N27697 10
D27697 N27697 0 diode
R27698 N27697 N27698 10
D27698 N27698 0 diode
R27699 N27698 N27699 10
D27699 N27699 0 diode
R27700 N27699 N27700 10
D27700 N27700 0 diode
R27701 N27700 N27701 10
D27701 N27701 0 diode
R27702 N27701 N27702 10
D27702 N27702 0 diode
R27703 N27702 N27703 10
D27703 N27703 0 diode
R27704 N27703 N27704 10
D27704 N27704 0 diode
R27705 N27704 N27705 10
D27705 N27705 0 diode
R27706 N27705 N27706 10
D27706 N27706 0 diode
R27707 N27706 N27707 10
D27707 N27707 0 diode
R27708 N27707 N27708 10
D27708 N27708 0 diode
R27709 N27708 N27709 10
D27709 N27709 0 diode
R27710 N27709 N27710 10
D27710 N27710 0 diode
R27711 N27710 N27711 10
D27711 N27711 0 diode
R27712 N27711 N27712 10
D27712 N27712 0 diode
R27713 N27712 N27713 10
D27713 N27713 0 diode
R27714 N27713 N27714 10
D27714 N27714 0 diode
R27715 N27714 N27715 10
D27715 N27715 0 diode
R27716 N27715 N27716 10
D27716 N27716 0 diode
R27717 N27716 N27717 10
D27717 N27717 0 diode
R27718 N27717 N27718 10
D27718 N27718 0 diode
R27719 N27718 N27719 10
D27719 N27719 0 diode
R27720 N27719 N27720 10
D27720 N27720 0 diode
R27721 N27720 N27721 10
D27721 N27721 0 diode
R27722 N27721 N27722 10
D27722 N27722 0 diode
R27723 N27722 N27723 10
D27723 N27723 0 diode
R27724 N27723 N27724 10
D27724 N27724 0 diode
R27725 N27724 N27725 10
D27725 N27725 0 diode
R27726 N27725 N27726 10
D27726 N27726 0 diode
R27727 N27726 N27727 10
D27727 N27727 0 diode
R27728 N27727 N27728 10
D27728 N27728 0 diode
R27729 N27728 N27729 10
D27729 N27729 0 diode
R27730 N27729 N27730 10
D27730 N27730 0 diode
R27731 N27730 N27731 10
D27731 N27731 0 diode
R27732 N27731 N27732 10
D27732 N27732 0 diode
R27733 N27732 N27733 10
D27733 N27733 0 diode
R27734 N27733 N27734 10
D27734 N27734 0 diode
R27735 N27734 N27735 10
D27735 N27735 0 diode
R27736 N27735 N27736 10
D27736 N27736 0 diode
R27737 N27736 N27737 10
D27737 N27737 0 diode
R27738 N27737 N27738 10
D27738 N27738 0 diode
R27739 N27738 N27739 10
D27739 N27739 0 diode
R27740 N27739 N27740 10
D27740 N27740 0 diode
R27741 N27740 N27741 10
D27741 N27741 0 diode
R27742 N27741 N27742 10
D27742 N27742 0 diode
R27743 N27742 N27743 10
D27743 N27743 0 diode
R27744 N27743 N27744 10
D27744 N27744 0 diode
R27745 N27744 N27745 10
D27745 N27745 0 diode
R27746 N27745 N27746 10
D27746 N27746 0 diode
R27747 N27746 N27747 10
D27747 N27747 0 diode
R27748 N27747 N27748 10
D27748 N27748 0 diode
R27749 N27748 N27749 10
D27749 N27749 0 diode
R27750 N27749 N27750 10
D27750 N27750 0 diode
R27751 N27750 N27751 10
D27751 N27751 0 diode
R27752 N27751 N27752 10
D27752 N27752 0 diode
R27753 N27752 N27753 10
D27753 N27753 0 diode
R27754 N27753 N27754 10
D27754 N27754 0 diode
R27755 N27754 N27755 10
D27755 N27755 0 diode
R27756 N27755 N27756 10
D27756 N27756 0 diode
R27757 N27756 N27757 10
D27757 N27757 0 diode
R27758 N27757 N27758 10
D27758 N27758 0 diode
R27759 N27758 N27759 10
D27759 N27759 0 diode
R27760 N27759 N27760 10
D27760 N27760 0 diode
R27761 N27760 N27761 10
D27761 N27761 0 diode
R27762 N27761 N27762 10
D27762 N27762 0 diode
R27763 N27762 N27763 10
D27763 N27763 0 diode
R27764 N27763 N27764 10
D27764 N27764 0 diode
R27765 N27764 N27765 10
D27765 N27765 0 diode
R27766 N27765 N27766 10
D27766 N27766 0 diode
R27767 N27766 N27767 10
D27767 N27767 0 diode
R27768 N27767 N27768 10
D27768 N27768 0 diode
R27769 N27768 N27769 10
D27769 N27769 0 diode
R27770 N27769 N27770 10
D27770 N27770 0 diode
R27771 N27770 N27771 10
D27771 N27771 0 diode
R27772 N27771 N27772 10
D27772 N27772 0 diode
R27773 N27772 N27773 10
D27773 N27773 0 diode
R27774 N27773 N27774 10
D27774 N27774 0 diode
R27775 N27774 N27775 10
D27775 N27775 0 diode
R27776 N27775 N27776 10
D27776 N27776 0 diode
R27777 N27776 N27777 10
D27777 N27777 0 diode
R27778 N27777 N27778 10
D27778 N27778 0 diode
R27779 N27778 N27779 10
D27779 N27779 0 diode
R27780 N27779 N27780 10
D27780 N27780 0 diode
R27781 N27780 N27781 10
D27781 N27781 0 diode
R27782 N27781 N27782 10
D27782 N27782 0 diode
R27783 N27782 N27783 10
D27783 N27783 0 diode
R27784 N27783 N27784 10
D27784 N27784 0 diode
R27785 N27784 N27785 10
D27785 N27785 0 diode
R27786 N27785 N27786 10
D27786 N27786 0 diode
R27787 N27786 N27787 10
D27787 N27787 0 diode
R27788 N27787 N27788 10
D27788 N27788 0 diode
R27789 N27788 N27789 10
D27789 N27789 0 diode
R27790 N27789 N27790 10
D27790 N27790 0 diode
R27791 N27790 N27791 10
D27791 N27791 0 diode
R27792 N27791 N27792 10
D27792 N27792 0 diode
R27793 N27792 N27793 10
D27793 N27793 0 diode
R27794 N27793 N27794 10
D27794 N27794 0 diode
R27795 N27794 N27795 10
D27795 N27795 0 diode
R27796 N27795 N27796 10
D27796 N27796 0 diode
R27797 N27796 N27797 10
D27797 N27797 0 diode
R27798 N27797 N27798 10
D27798 N27798 0 diode
R27799 N27798 N27799 10
D27799 N27799 0 diode
R27800 N27799 N27800 10
D27800 N27800 0 diode
R27801 N27800 N27801 10
D27801 N27801 0 diode
R27802 N27801 N27802 10
D27802 N27802 0 diode
R27803 N27802 N27803 10
D27803 N27803 0 diode
R27804 N27803 N27804 10
D27804 N27804 0 diode
R27805 N27804 N27805 10
D27805 N27805 0 diode
R27806 N27805 N27806 10
D27806 N27806 0 diode
R27807 N27806 N27807 10
D27807 N27807 0 diode
R27808 N27807 N27808 10
D27808 N27808 0 diode
R27809 N27808 N27809 10
D27809 N27809 0 diode
R27810 N27809 N27810 10
D27810 N27810 0 diode
R27811 N27810 N27811 10
D27811 N27811 0 diode
R27812 N27811 N27812 10
D27812 N27812 0 diode
R27813 N27812 N27813 10
D27813 N27813 0 diode
R27814 N27813 N27814 10
D27814 N27814 0 diode
R27815 N27814 N27815 10
D27815 N27815 0 diode
R27816 N27815 N27816 10
D27816 N27816 0 diode
R27817 N27816 N27817 10
D27817 N27817 0 diode
R27818 N27817 N27818 10
D27818 N27818 0 diode
R27819 N27818 N27819 10
D27819 N27819 0 diode
R27820 N27819 N27820 10
D27820 N27820 0 diode
R27821 N27820 N27821 10
D27821 N27821 0 diode
R27822 N27821 N27822 10
D27822 N27822 0 diode
R27823 N27822 N27823 10
D27823 N27823 0 diode
R27824 N27823 N27824 10
D27824 N27824 0 diode
R27825 N27824 N27825 10
D27825 N27825 0 diode
R27826 N27825 N27826 10
D27826 N27826 0 diode
R27827 N27826 N27827 10
D27827 N27827 0 diode
R27828 N27827 N27828 10
D27828 N27828 0 diode
R27829 N27828 N27829 10
D27829 N27829 0 diode
R27830 N27829 N27830 10
D27830 N27830 0 diode
R27831 N27830 N27831 10
D27831 N27831 0 diode
R27832 N27831 N27832 10
D27832 N27832 0 diode
R27833 N27832 N27833 10
D27833 N27833 0 diode
R27834 N27833 N27834 10
D27834 N27834 0 diode
R27835 N27834 N27835 10
D27835 N27835 0 diode
R27836 N27835 N27836 10
D27836 N27836 0 diode
R27837 N27836 N27837 10
D27837 N27837 0 diode
R27838 N27837 N27838 10
D27838 N27838 0 diode
R27839 N27838 N27839 10
D27839 N27839 0 diode
R27840 N27839 N27840 10
D27840 N27840 0 diode
R27841 N27840 N27841 10
D27841 N27841 0 diode
R27842 N27841 N27842 10
D27842 N27842 0 diode
R27843 N27842 N27843 10
D27843 N27843 0 diode
R27844 N27843 N27844 10
D27844 N27844 0 diode
R27845 N27844 N27845 10
D27845 N27845 0 diode
R27846 N27845 N27846 10
D27846 N27846 0 diode
R27847 N27846 N27847 10
D27847 N27847 0 diode
R27848 N27847 N27848 10
D27848 N27848 0 diode
R27849 N27848 N27849 10
D27849 N27849 0 diode
R27850 N27849 N27850 10
D27850 N27850 0 diode
R27851 N27850 N27851 10
D27851 N27851 0 diode
R27852 N27851 N27852 10
D27852 N27852 0 diode
R27853 N27852 N27853 10
D27853 N27853 0 diode
R27854 N27853 N27854 10
D27854 N27854 0 diode
R27855 N27854 N27855 10
D27855 N27855 0 diode
R27856 N27855 N27856 10
D27856 N27856 0 diode
R27857 N27856 N27857 10
D27857 N27857 0 diode
R27858 N27857 N27858 10
D27858 N27858 0 diode
R27859 N27858 N27859 10
D27859 N27859 0 diode
R27860 N27859 N27860 10
D27860 N27860 0 diode
R27861 N27860 N27861 10
D27861 N27861 0 diode
R27862 N27861 N27862 10
D27862 N27862 0 diode
R27863 N27862 N27863 10
D27863 N27863 0 diode
R27864 N27863 N27864 10
D27864 N27864 0 diode
R27865 N27864 N27865 10
D27865 N27865 0 diode
R27866 N27865 N27866 10
D27866 N27866 0 diode
R27867 N27866 N27867 10
D27867 N27867 0 diode
R27868 N27867 N27868 10
D27868 N27868 0 diode
R27869 N27868 N27869 10
D27869 N27869 0 diode
R27870 N27869 N27870 10
D27870 N27870 0 diode
R27871 N27870 N27871 10
D27871 N27871 0 diode
R27872 N27871 N27872 10
D27872 N27872 0 diode
R27873 N27872 N27873 10
D27873 N27873 0 diode
R27874 N27873 N27874 10
D27874 N27874 0 diode
R27875 N27874 N27875 10
D27875 N27875 0 diode
R27876 N27875 N27876 10
D27876 N27876 0 diode
R27877 N27876 N27877 10
D27877 N27877 0 diode
R27878 N27877 N27878 10
D27878 N27878 0 diode
R27879 N27878 N27879 10
D27879 N27879 0 diode
R27880 N27879 N27880 10
D27880 N27880 0 diode
R27881 N27880 N27881 10
D27881 N27881 0 diode
R27882 N27881 N27882 10
D27882 N27882 0 diode
R27883 N27882 N27883 10
D27883 N27883 0 diode
R27884 N27883 N27884 10
D27884 N27884 0 diode
R27885 N27884 N27885 10
D27885 N27885 0 diode
R27886 N27885 N27886 10
D27886 N27886 0 diode
R27887 N27886 N27887 10
D27887 N27887 0 diode
R27888 N27887 N27888 10
D27888 N27888 0 diode
R27889 N27888 N27889 10
D27889 N27889 0 diode
R27890 N27889 N27890 10
D27890 N27890 0 diode
R27891 N27890 N27891 10
D27891 N27891 0 diode
R27892 N27891 N27892 10
D27892 N27892 0 diode
R27893 N27892 N27893 10
D27893 N27893 0 diode
R27894 N27893 N27894 10
D27894 N27894 0 diode
R27895 N27894 N27895 10
D27895 N27895 0 diode
R27896 N27895 N27896 10
D27896 N27896 0 diode
R27897 N27896 N27897 10
D27897 N27897 0 diode
R27898 N27897 N27898 10
D27898 N27898 0 diode
R27899 N27898 N27899 10
D27899 N27899 0 diode
R27900 N27899 N27900 10
D27900 N27900 0 diode
R27901 N27900 N27901 10
D27901 N27901 0 diode
R27902 N27901 N27902 10
D27902 N27902 0 diode
R27903 N27902 N27903 10
D27903 N27903 0 diode
R27904 N27903 N27904 10
D27904 N27904 0 diode
R27905 N27904 N27905 10
D27905 N27905 0 diode
R27906 N27905 N27906 10
D27906 N27906 0 diode
R27907 N27906 N27907 10
D27907 N27907 0 diode
R27908 N27907 N27908 10
D27908 N27908 0 diode
R27909 N27908 N27909 10
D27909 N27909 0 diode
R27910 N27909 N27910 10
D27910 N27910 0 diode
R27911 N27910 N27911 10
D27911 N27911 0 diode
R27912 N27911 N27912 10
D27912 N27912 0 diode
R27913 N27912 N27913 10
D27913 N27913 0 diode
R27914 N27913 N27914 10
D27914 N27914 0 diode
R27915 N27914 N27915 10
D27915 N27915 0 diode
R27916 N27915 N27916 10
D27916 N27916 0 diode
R27917 N27916 N27917 10
D27917 N27917 0 diode
R27918 N27917 N27918 10
D27918 N27918 0 diode
R27919 N27918 N27919 10
D27919 N27919 0 diode
R27920 N27919 N27920 10
D27920 N27920 0 diode
R27921 N27920 N27921 10
D27921 N27921 0 diode
R27922 N27921 N27922 10
D27922 N27922 0 diode
R27923 N27922 N27923 10
D27923 N27923 0 diode
R27924 N27923 N27924 10
D27924 N27924 0 diode
R27925 N27924 N27925 10
D27925 N27925 0 diode
R27926 N27925 N27926 10
D27926 N27926 0 diode
R27927 N27926 N27927 10
D27927 N27927 0 diode
R27928 N27927 N27928 10
D27928 N27928 0 diode
R27929 N27928 N27929 10
D27929 N27929 0 diode
R27930 N27929 N27930 10
D27930 N27930 0 diode
R27931 N27930 N27931 10
D27931 N27931 0 diode
R27932 N27931 N27932 10
D27932 N27932 0 diode
R27933 N27932 N27933 10
D27933 N27933 0 diode
R27934 N27933 N27934 10
D27934 N27934 0 diode
R27935 N27934 N27935 10
D27935 N27935 0 diode
R27936 N27935 N27936 10
D27936 N27936 0 diode
R27937 N27936 N27937 10
D27937 N27937 0 diode
R27938 N27937 N27938 10
D27938 N27938 0 diode
R27939 N27938 N27939 10
D27939 N27939 0 diode
R27940 N27939 N27940 10
D27940 N27940 0 diode
R27941 N27940 N27941 10
D27941 N27941 0 diode
R27942 N27941 N27942 10
D27942 N27942 0 diode
R27943 N27942 N27943 10
D27943 N27943 0 diode
R27944 N27943 N27944 10
D27944 N27944 0 diode
R27945 N27944 N27945 10
D27945 N27945 0 diode
R27946 N27945 N27946 10
D27946 N27946 0 diode
R27947 N27946 N27947 10
D27947 N27947 0 diode
R27948 N27947 N27948 10
D27948 N27948 0 diode
R27949 N27948 N27949 10
D27949 N27949 0 diode
R27950 N27949 N27950 10
D27950 N27950 0 diode
R27951 N27950 N27951 10
D27951 N27951 0 diode
R27952 N27951 N27952 10
D27952 N27952 0 diode
R27953 N27952 N27953 10
D27953 N27953 0 diode
R27954 N27953 N27954 10
D27954 N27954 0 diode
R27955 N27954 N27955 10
D27955 N27955 0 diode
R27956 N27955 N27956 10
D27956 N27956 0 diode
R27957 N27956 N27957 10
D27957 N27957 0 diode
R27958 N27957 N27958 10
D27958 N27958 0 diode
R27959 N27958 N27959 10
D27959 N27959 0 diode
R27960 N27959 N27960 10
D27960 N27960 0 diode
R27961 N27960 N27961 10
D27961 N27961 0 diode
R27962 N27961 N27962 10
D27962 N27962 0 diode
R27963 N27962 N27963 10
D27963 N27963 0 diode
R27964 N27963 N27964 10
D27964 N27964 0 diode
R27965 N27964 N27965 10
D27965 N27965 0 diode
R27966 N27965 N27966 10
D27966 N27966 0 diode
R27967 N27966 N27967 10
D27967 N27967 0 diode
R27968 N27967 N27968 10
D27968 N27968 0 diode
R27969 N27968 N27969 10
D27969 N27969 0 diode
R27970 N27969 N27970 10
D27970 N27970 0 diode
R27971 N27970 N27971 10
D27971 N27971 0 diode
R27972 N27971 N27972 10
D27972 N27972 0 diode
R27973 N27972 N27973 10
D27973 N27973 0 diode
R27974 N27973 N27974 10
D27974 N27974 0 diode
R27975 N27974 N27975 10
D27975 N27975 0 diode
R27976 N27975 N27976 10
D27976 N27976 0 diode
R27977 N27976 N27977 10
D27977 N27977 0 diode
R27978 N27977 N27978 10
D27978 N27978 0 diode
R27979 N27978 N27979 10
D27979 N27979 0 diode
R27980 N27979 N27980 10
D27980 N27980 0 diode
R27981 N27980 N27981 10
D27981 N27981 0 diode
R27982 N27981 N27982 10
D27982 N27982 0 diode
R27983 N27982 N27983 10
D27983 N27983 0 diode
R27984 N27983 N27984 10
D27984 N27984 0 diode
R27985 N27984 N27985 10
D27985 N27985 0 diode
R27986 N27985 N27986 10
D27986 N27986 0 diode
R27987 N27986 N27987 10
D27987 N27987 0 diode
R27988 N27987 N27988 10
D27988 N27988 0 diode
R27989 N27988 N27989 10
D27989 N27989 0 diode
R27990 N27989 N27990 10
D27990 N27990 0 diode
R27991 N27990 N27991 10
D27991 N27991 0 diode
R27992 N27991 N27992 10
D27992 N27992 0 diode
R27993 N27992 N27993 10
D27993 N27993 0 diode
R27994 N27993 N27994 10
D27994 N27994 0 diode
R27995 N27994 N27995 10
D27995 N27995 0 diode
R27996 N27995 N27996 10
D27996 N27996 0 diode
R27997 N27996 N27997 10
D27997 N27997 0 diode
R27998 N27997 N27998 10
D27998 N27998 0 diode
R27999 N27998 N27999 10
D27999 N27999 0 diode
R28000 N27999 N28000 10
D28000 N28000 0 diode
R28001 N28000 N28001 10
D28001 N28001 0 diode
R28002 N28001 N28002 10
D28002 N28002 0 diode
R28003 N28002 N28003 10
D28003 N28003 0 diode
R28004 N28003 N28004 10
D28004 N28004 0 diode
R28005 N28004 N28005 10
D28005 N28005 0 diode
R28006 N28005 N28006 10
D28006 N28006 0 diode
R28007 N28006 N28007 10
D28007 N28007 0 diode
R28008 N28007 N28008 10
D28008 N28008 0 diode
R28009 N28008 N28009 10
D28009 N28009 0 diode
R28010 N28009 N28010 10
D28010 N28010 0 diode
R28011 N28010 N28011 10
D28011 N28011 0 diode
R28012 N28011 N28012 10
D28012 N28012 0 diode
R28013 N28012 N28013 10
D28013 N28013 0 diode
R28014 N28013 N28014 10
D28014 N28014 0 diode
R28015 N28014 N28015 10
D28015 N28015 0 diode
R28016 N28015 N28016 10
D28016 N28016 0 diode
R28017 N28016 N28017 10
D28017 N28017 0 diode
R28018 N28017 N28018 10
D28018 N28018 0 diode
R28019 N28018 N28019 10
D28019 N28019 0 diode
R28020 N28019 N28020 10
D28020 N28020 0 diode
R28021 N28020 N28021 10
D28021 N28021 0 diode
R28022 N28021 N28022 10
D28022 N28022 0 diode
R28023 N28022 N28023 10
D28023 N28023 0 diode
R28024 N28023 N28024 10
D28024 N28024 0 diode
R28025 N28024 N28025 10
D28025 N28025 0 diode
R28026 N28025 N28026 10
D28026 N28026 0 diode
R28027 N28026 N28027 10
D28027 N28027 0 diode
R28028 N28027 N28028 10
D28028 N28028 0 diode
R28029 N28028 N28029 10
D28029 N28029 0 diode
R28030 N28029 N28030 10
D28030 N28030 0 diode
R28031 N28030 N28031 10
D28031 N28031 0 diode
R28032 N28031 N28032 10
D28032 N28032 0 diode
R28033 N28032 N28033 10
D28033 N28033 0 diode
R28034 N28033 N28034 10
D28034 N28034 0 diode
R28035 N28034 N28035 10
D28035 N28035 0 diode
R28036 N28035 N28036 10
D28036 N28036 0 diode
R28037 N28036 N28037 10
D28037 N28037 0 diode
R28038 N28037 N28038 10
D28038 N28038 0 diode
R28039 N28038 N28039 10
D28039 N28039 0 diode
R28040 N28039 N28040 10
D28040 N28040 0 diode
R28041 N28040 N28041 10
D28041 N28041 0 diode
R28042 N28041 N28042 10
D28042 N28042 0 diode
R28043 N28042 N28043 10
D28043 N28043 0 diode
R28044 N28043 N28044 10
D28044 N28044 0 diode
R28045 N28044 N28045 10
D28045 N28045 0 diode
R28046 N28045 N28046 10
D28046 N28046 0 diode
R28047 N28046 N28047 10
D28047 N28047 0 diode
R28048 N28047 N28048 10
D28048 N28048 0 diode
R28049 N28048 N28049 10
D28049 N28049 0 diode
R28050 N28049 N28050 10
D28050 N28050 0 diode
R28051 N28050 N28051 10
D28051 N28051 0 diode
R28052 N28051 N28052 10
D28052 N28052 0 diode
R28053 N28052 N28053 10
D28053 N28053 0 diode
R28054 N28053 N28054 10
D28054 N28054 0 diode
R28055 N28054 N28055 10
D28055 N28055 0 diode
R28056 N28055 N28056 10
D28056 N28056 0 diode
R28057 N28056 N28057 10
D28057 N28057 0 diode
R28058 N28057 N28058 10
D28058 N28058 0 diode
R28059 N28058 N28059 10
D28059 N28059 0 diode
R28060 N28059 N28060 10
D28060 N28060 0 diode
R28061 N28060 N28061 10
D28061 N28061 0 diode
R28062 N28061 N28062 10
D28062 N28062 0 diode
R28063 N28062 N28063 10
D28063 N28063 0 diode
R28064 N28063 N28064 10
D28064 N28064 0 diode
R28065 N28064 N28065 10
D28065 N28065 0 diode
R28066 N28065 N28066 10
D28066 N28066 0 diode
R28067 N28066 N28067 10
D28067 N28067 0 diode
R28068 N28067 N28068 10
D28068 N28068 0 diode
R28069 N28068 N28069 10
D28069 N28069 0 diode
R28070 N28069 N28070 10
D28070 N28070 0 diode
R28071 N28070 N28071 10
D28071 N28071 0 diode
R28072 N28071 N28072 10
D28072 N28072 0 diode
R28073 N28072 N28073 10
D28073 N28073 0 diode
R28074 N28073 N28074 10
D28074 N28074 0 diode
R28075 N28074 N28075 10
D28075 N28075 0 diode
R28076 N28075 N28076 10
D28076 N28076 0 diode
R28077 N28076 N28077 10
D28077 N28077 0 diode
R28078 N28077 N28078 10
D28078 N28078 0 diode
R28079 N28078 N28079 10
D28079 N28079 0 diode
R28080 N28079 N28080 10
D28080 N28080 0 diode
R28081 N28080 N28081 10
D28081 N28081 0 diode
R28082 N28081 N28082 10
D28082 N28082 0 diode
R28083 N28082 N28083 10
D28083 N28083 0 diode
R28084 N28083 N28084 10
D28084 N28084 0 diode
R28085 N28084 N28085 10
D28085 N28085 0 diode
R28086 N28085 N28086 10
D28086 N28086 0 diode
R28087 N28086 N28087 10
D28087 N28087 0 diode
R28088 N28087 N28088 10
D28088 N28088 0 diode
R28089 N28088 N28089 10
D28089 N28089 0 diode
R28090 N28089 N28090 10
D28090 N28090 0 diode
R28091 N28090 N28091 10
D28091 N28091 0 diode
R28092 N28091 N28092 10
D28092 N28092 0 diode
R28093 N28092 N28093 10
D28093 N28093 0 diode
R28094 N28093 N28094 10
D28094 N28094 0 diode
R28095 N28094 N28095 10
D28095 N28095 0 diode
R28096 N28095 N28096 10
D28096 N28096 0 diode
R28097 N28096 N28097 10
D28097 N28097 0 diode
R28098 N28097 N28098 10
D28098 N28098 0 diode
R28099 N28098 N28099 10
D28099 N28099 0 diode
R28100 N28099 N28100 10
D28100 N28100 0 diode
R28101 N28100 N28101 10
D28101 N28101 0 diode
R28102 N28101 N28102 10
D28102 N28102 0 diode
R28103 N28102 N28103 10
D28103 N28103 0 diode
R28104 N28103 N28104 10
D28104 N28104 0 diode
R28105 N28104 N28105 10
D28105 N28105 0 diode
R28106 N28105 N28106 10
D28106 N28106 0 diode
R28107 N28106 N28107 10
D28107 N28107 0 diode
R28108 N28107 N28108 10
D28108 N28108 0 diode
R28109 N28108 N28109 10
D28109 N28109 0 diode
R28110 N28109 N28110 10
D28110 N28110 0 diode
R28111 N28110 N28111 10
D28111 N28111 0 diode
R28112 N28111 N28112 10
D28112 N28112 0 diode
R28113 N28112 N28113 10
D28113 N28113 0 diode
R28114 N28113 N28114 10
D28114 N28114 0 diode
R28115 N28114 N28115 10
D28115 N28115 0 diode
R28116 N28115 N28116 10
D28116 N28116 0 diode
R28117 N28116 N28117 10
D28117 N28117 0 diode
R28118 N28117 N28118 10
D28118 N28118 0 diode
R28119 N28118 N28119 10
D28119 N28119 0 diode
R28120 N28119 N28120 10
D28120 N28120 0 diode
R28121 N28120 N28121 10
D28121 N28121 0 diode
R28122 N28121 N28122 10
D28122 N28122 0 diode
R28123 N28122 N28123 10
D28123 N28123 0 diode
R28124 N28123 N28124 10
D28124 N28124 0 diode
R28125 N28124 N28125 10
D28125 N28125 0 diode
R28126 N28125 N28126 10
D28126 N28126 0 diode
R28127 N28126 N28127 10
D28127 N28127 0 diode
R28128 N28127 N28128 10
D28128 N28128 0 diode
R28129 N28128 N28129 10
D28129 N28129 0 diode
R28130 N28129 N28130 10
D28130 N28130 0 diode
R28131 N28130 N28131 10
D28131 N28131 0 diode
R28132 N28131 N28132 10
D28132 N28132 0 diode
R28133 N28132 N28133 10
D28133 N28133 0 diode
R28134 N28133 N28134 10
D28134 N28134 0 diode
R28135 N28134 N28135 10
D28135 N28135 0 diode
R28136 N28135 N28136 10
D28136 N28136 0 diode
R28137 N28136 N28137 10
D28137 N28137 0 diode
R28138 N28137 N28138 10
D28138 N28138 0 diode
R28139 N28138 N28139 10
D28139 N28139 0 diode
R28140 N28139 N28140 10
D28140 N28140 0 diode
R28141 N28140 N28141 10
D28141 N28141 0 diode
R28142 N28141 N28142 10
D28142 N28142 0 diode
R28143 N28142 N28143 10
D28143 N28143 0 diode
R28144 N28143 N28144 10
D28144 N28144 0 diode
R28145 N28144 N28145 10
D28145 N28145 0 diode
R28146 N28145 N28146 10
D28146 N28146 0 diode
R28147 N28146 N28147 10
D28147 N28147 0 diode
R28148 N28147 N28148 10
D28148 N28148 0 diode
R28149 N28148 N28149 10
D28149 N28149 0 diode
R28150 N28149 N28150 10
D28150 N28150 0 diode
R28151 N28150 N28151 10
D28151 N28151 0 diode
R28152 N28151 N28152 10
D28152 N28152 0 diode
R28153 N28152 N28153 10
D28153 N28153 0 diode
R28154 N28153 N28154 10
D28154 N28154 0 diode
R28155 N28154 N28155 10
D28155 N28155 0 diode
R28156 N28155 N28156 10
D28156 N28156 0 diode
R28157 N28156 N28157 10
D28157 N28157 0 diode
R28158 N28157 N28158 10
D28158 N28158 0 diode
R28159 N28158 N28159 10
D28159 N28159 0 diode
R28160 N28159 N28160 10
D28160 N28160 0 diode
R28161 N28160 N28161 10
D28161 N28161 0 diode
R28162 N28161 N28162 10
D28162 N28162 0 diode
R28163 N28162 N28163 10
D28163 N28163 0 diode
R28164 N28163 N28164 10
D28164 N28164 0 diode
R28165 N28164 N28165 10
D28165 N28165 0 diode
R28166 N28165 N28166 10
D28166 N28166 0 diode
R28167 N28166 N28167 10
D28167 N28167 0 diode
R28168 N28167 N28168 10
D28168 N28168 0 diode
R28169 N28168 N28169 10
D28169 N28169 0 diode
R28170 N28169 N28170 10
D28170 N28170 0 diode
R28171 N28170 N28171 10
D28171 N28171 0 diode
R28172 N28171 N28172 10
D28172 N28172 0 diode
R28173 N28172 N28173 10
D28173 N28173 0 diode
R28174 N28173 N28174 10
D28174 N28174 0 diode
R28175 N28174 N28175 10
D28175 N28175 0 diode
R28176 N28175 N28176 10
D28176 N28176 0 diode
R28177 N28176 N28177 10
D28177 N28177 0 diode
R28178 N28177 N28178 10
D28178 N28178 0 diode
R28179 N28178 N28179 10
D28179 N28179 0 diode
R28180 N28179 N28180 10
D28180 N28180 0 diode
R28181 N28180 N28181 10
D28181 N28181 0 diode
R28182 N28181 N28182 10
D28182 N28182 0 diode
R28183 N28182 N28183 10
D28183 N28183 0 diode
R28184 N28183 N28184 10
D28184 N28184 0 diode
R28185 N28184 N28185 10
D28185 N28185 0 diode
R28186 N28185 N28186 10
D28186 N28186 0 diode
R28187 N28186 N28187 10
D28187 N28187 0 diode
R28188 N28187 N28188 10
D28188 N28188 0 diode
R28189 N28188 N28189 10
D28189 N28189 0 diode
R28190 N28189 N28190 10
D28190 N28190 0 diode
R28191 N28190 N28191 10
D28191 N28191 0 diode
R28192 N28191 N28192 10
D28192 N28192 0 diode
R28193 N28192 N28193 10
D28193 N28193 0 diode
R28194 N28193 N28194 10
D28194 N28194 0 diode
R28195 N28194 N28195 10
D28195 N28195 0 diode
R28196 N28195 N28196 10
D28196 N28196 0 diode
R28197 N28196 N28197 10
D28197 N28197 0 diode
R28198 N28197 N28198 10
D28198 N28198 0 diode
R28199 N28198 N28199 10
D28199 N28199 0 diode
R28200 N28199 N28200 10
D28200 N28200 0 diode
R28201 N28200 N28201 10
D28201 N28201 0 diode
R28202 N28201 N28202 10
D28202 N28202 0 diode
R28203 N28202 N28203 10
D28203 N28203 0 diode
R28204 N28203 N28204 10
D28204 N28204 0 diode
R28205 N28204 N28205 10
D28205 N28205 0 diode
R28206 N28205 N28206 10
D28206 N28206 0 diode
R28207 N28206 N28207 10
D28207 N28207 0 diode
R28208 N28207 N28208 10
D28208 N28208 0 diode
R28209 N28208 N28209 10
D28209 N28209 0 diode
R28210 N28209 N28210 10
D28210 N28210 0 diode
R28211 N28210 N28211 10
D28211 N28211 0 diode
R28212 N28211 N28212 10
D28212 N28212 0 diode
R28213 N28212 N28213 10
D28213 N28213 0 diode
R28214 N28213 N28214 10
D28214 N28214 0 diode
R28215 N28214 N28215 10
D28215 N28215 0 diode
R28216 N28215 N28216 10
D28216 N28216 0 diode
R28217 N28216 N28217 10
D28217 N28217 0 diode
R28218 N28217 N28218 10
D28218 N28218 0 diode
R28219 N28218 N28219 10
D28219 N28219 0 diode
R28220 N28219 N28220 10
D28220 N28220 0 diode
R28221 N28220 N28221 10
D28221 N28221 0 diode
R28222 N28221 N28222 10
D28222 N28222 0 diode
R28223 N28222 N28223 10
D28223 N28223 0 diode
R28224 N28223 N28224 10
D28224 N28224 0 diode
R28225 N28224 N28225 10
D28225 N28225 0 diode
R28226 N28225 N28226 10
D28226 N28226 0 diode
R28227 N28226 N28227 10
D28227 N28227 0 diode
R28228 N28227 N28228 10
D28228 N28228 0 diode
R28229 N28228 N28229 10
D28229 N28229 0 diode
R28230 N28229 N28230 10
D28230 N28230 0 diode
R28231 N28230 N28231 10
D28231 N28231 0 diode
R28232 N28231 N28232 10
D28232 N28232 0 diode
R28233 N28232 N28233 10
D28233 N28233 0 diode
R28234 N28233 N28234 10
D28234 N28234 0 diode
R28235 N28234 N28235 10
D28235 N28235 0 diode
R28236 N28235 N28236 10
D28236 N28236 0 diode
R28237 N28236 N28237 10
D28237 N28237 0 diode
R28238 N28237 N28238 10
D28238 N28238 0 diode
R28239 N28238 N28239 10
D28239 N28239 0 diode
R28240 N28239 N28240 10
D28240 N28240 0 diode
R28241 N28240 N28241 10
D28241 N28241 0 diode
R28242 N28241 N28242 10
D28242 N28242 0 diode
R28243 N28242 N28243 10
D28243 N28243 0 diode
R28244 N28243 N28244 10
D28244 N28244 0 diode
R28245 N28244 N28245 10
D28245 N28245 0 diode
R28246 N28245 N28246 10
D28246 N28246 0 diode
R28247 N28246 N28247 10
D28247 N28247 0 diode
R28248 N28247 N28248 10
D28248 N28248 0 diode
R28249 N28248 N28249 10
D28249 N28249 0 diode
R28250 N28249 N28250 10
D28250 N28250 0 diode
R28251 N28250 N28251 10
D28251 N28251 0 diode
R28252 N28251 N28252 10
D28252 N28252 0 diode
R28253 N28252 N28253 10
D28253 N28253 0 diode
R28254 N28253 N28254 10
D28254 N28254 0 diode
R28255 N28254 N28255 10
D28255 N28255 0 diode
R28256 N28255 N28256 10
D28256 N28256 0 diode
R28257 N28256 N28257 10
D28257 N28257 0 diode
R28258 N28257 N28258 10
D28258 N28258 0 diode
R28259 N28258 N28259 10
D28259 N28259 0 diode
R28260 N28259 N28260 10
D28260 N28260 0 diode
R28261 N28260 N28261 10
D28261 N28261 0 diode
R28262 N28261 N28262 10
D28262 N28262 0 diode
R28263 N28262 N28263 10
D28263 N28263 0 diode
R28264 N28263 N28264 10
D28264 N28264 0 diode
R28265 N28264 N28265 10
D28265 N28265 0 diode
R28266 N28265 N28266 10
D28266 N28266 0 diode
R28267 N28266 N28267 10
D28267 N28267 0 diode
R28268 N28267 N28268 10
D28268 N28268 0 diode
R28269 N28268 N28269 10
D28269 N28269 0 diode
R28270 N28269 N28270 10
D28270 N28270 0 diode
R28271 N28270 N28271 10
D28271 N28271 0 diode
R28272 N28271 N28272 10
D28272 N28272 0 diode
R28273 N28272 N28273 10
D28273 N28273 0 diode
R28274 N28273 N28274 10
D28274 N28274 0 diode
R28275 N28274 N28275 10
D28275 N28275 0 diode
R28276 N28275 N28276 10
D28276 N28276 0 diode
R28277 N28276 N28277 10
D28277 N28277 0 diode
R28278 N28277 N28278 10
D28278 N28278 0 diode
R28279 N28278 N28279 10
D28279 N28279 0 diode
R28280 N28279 N28280 10
D28280 N28280 0 diode
R28281 N28280 N28281 10
D28281 N28281 0 diode
R28282 N28281 N28282 10
D28282 N28282 0 diode
R28283 N28282 N28283 10
D28283 N28283 0 diode
R28284 N28283 N28284 10
D28284 N28284 0 diode
R28285 N28284 N28285 10
D28285 N28285 0 diode
R28286 N28285 N28286 10
D28286 N28286 0 diode
R28287 N28286 N28287 10
D28287 N28287 0 diode
R28288 N28287 N28288 10
D28288 N28288 0 diode
R28289 N28288 N28289 10
D28289 N28289 0 diode
R28290 N28289 N28290 10
D28290 N28290 0 diode
R28291 N28290 N28291 10
D28291 N28291 0 diode
R28292 N28291 N28292 10
D28292 N28292 0 diode
R28293 N28292 N28293 10
D28293 N28293 0 diode
R28294 N28293 N28294 10
D28294 N28294 0 diode
R28295 N28294 N28295 10
D28295 N28295 0 diode
R28296 N28295 N28296 10
D28296 N28296 0 diode
R28297 N28296 N28297 10
D28297 N28297 0 diode
R28298 N28297 N28298 10
D28298 N28298 0 diode
R28299 N28298 N28299 10
D28299 N28299 0 diode
R28300 N28299 N28300 10
D28300 N28300 0 diode
R28301 N28300 N28301 10
D28301 N28301 0 diode
R28302 N28301 N28302 10
D28302 N28302 0 diode
R28303 N28302 N28303 10
D28303 N28303 0 diode
R28304 N28303 N28304 10
D28304 N28304 0 diode
R28305 N28304 N28305 10
D28305 N28305 0 diode
R28306 N28305 N28306 10
D28306 N28306 0 diode
R28307 N28306 N28307 10
D28307 N28307 0 diode
R28308 N28307 N28308 10
D28308 N28308 0 diode
R28309 N28308 N28309 10
D28309 N28309 0 diode
R28310 N28309 N28310 10
D28310 N28310 0 diode
R28311 N28310 N28311 10
D28311 N28311 0 diode
R28312 N28311 N28312 10
D28312 N28312 0 diode
R28313 N28312 N28313 10
D28313 N28313 0 diode
R28314 N28313 N28314 10
D28314 N28314 0 diode
R28315 N28314 N28315 10
D28315 N28315 0 diode
R28316 N28315 N28316 10
D28316 N28316 0 diode
R28317 N28316 N28317 10
D28317 N28317 0 diode
R28318 N28317 N28318 10
D28318 N28318 0 diode
R28319 N28318 N28319 10
D28319 N28319 0 diode
R28320 N28319 N28320 10
D28320 N28320 0 diode
R28321 N28320 N28321 10
D28321 N28321 0 diode
R28322 N28321 N28322 10
D28322 N28322 0 diode
R28323 N28322 N28323 10
D28323 N28323 0 diode
R28324 N28323 N28324 10
D28324 N28324 0 diode
R28325 N28324 N28325 10
D28325 N28325 0 diode
R28326 N28325 N28326 10
D28326 N28326 0 diode
R28327 N28326 N28327 10
D28327 N28327 0 diode
R28328 N28327 N28328 10
D28328 N28328 0 diode
R28329 N28328 N28329 10
D28329 N28329 0 diode
R28330 N28329 N28330 10
D28330 N28330 0 diode
R28331 N28330 N28331 10
D28331 N28331 0 diode
R28332 N28331 N28332 10
D28332 N28332 0 diode
R28333 N28332 N28333 10
D28333 N28333 0 diode
R28334 N28333 N28334 10
D28334 N28334 0 diode
R28335 N28334 N28335 10
D28335 N28335 0 diode
R28336 N28335 N28336 10
D28336 N28336 0 diode
R28337 N28336 N28337 10
D28337 N28337 0 diode
R28338 N28337 N28338 10
D28338 N28338 0 diode
R28339 N28338 N28339 10
D28339 N28339 0 diode
R28340 N28339 N28340 10
D28340 N28340 0 diode
R28341 N28340 N28341 10
D28341 N28341 0 diode
R28342 N28341 N28342 10
D28342 N28342 0 diode
R28343 N28342 N28343 10
D28343 N28343 0 diode
R28344 N28343 N28344 10
D28344 N28344 0 diode
R28345 N28344 N28345 10
D28345 N28345 0 diode
R28346 N28345 N28346 10
D28346 N28346 0 diode
R28347 N28346 N28347 10
D28347 N28347 0 diode
R28348 N28347 N28348 10
D28348 N28348 0 diode
R28349 N28348 N28349 10
D28349 N28349 0 diode
R28350 N28349 N28350 10
D28350 N28350 0 diode
R28351 N28350 N28351 10
D28351 N28351 0 diode
R28352 N28351 N28352 10
D28352 N28352 0 diode
R28353 N28352 N28353 10
D28353 N28353 0 diode
R28354 N28353 N28354 10
D28354 N28354 0 diode
R28355 N28354 N28355 10
D28355 N28355 0 diode
R28356 N28355 N28356 10
D28356 N28356 0 diode
R28357 N28356 N28357 10
D28357 N28357 0 diode
R28358 N28357 N28358 10
D28358 N28358 0 diode
R28359 N28358 N28359 10
D28359 N28359 0 diode
R28360 N28359 N28360 10
D28360 N28360 0 diode
R28361 N28360 N28361 10
D28361 N28361 0 diode
R28362 N28361 N28362 10
D28362 N28362 0 diode
R28363 N28362 N28363 10
D28363 N28363 0 diode
R28364 N28363 N28364 10
D28364 N28364 0 diode
R28365 N28364 N28365 10
D28365 N28365 0 diode
R28366 N28365 N28366 10
D28366 N28366 0 diode
R28367 N28366 N28367 10
D28367 N28367 0 diode
R28368 N28367 N28368 10
D28368 N28368 0 diode
R28369 N28368 N28369 10
D28369 N28369 0 diode
R28370 N28369 N28370 10
D28370 N28370 0 diode
R28371 N28370 N28371 10
D28371 N28371 0 diode
R28372 N28371 N28372 10
D28372 N28372 0 diode
R28373 N28372 N28373 10
D28373 N28373 0 diode
R28374 N28373 N28374 10
D28374 N28374 0 diode
R28375 N28374 N28375 10
D28375 N28375 0 diode
R28376 N28375 N28376 10
D28376 N28376 0 diode
R28377 N28376 N28377 10
D28377 N28377 0 diode
R28378 N28377 N28378 10
D28378 N28378 0 diode
R28379 N28378 N28379 10
D28379 N28379 0 diode
R28380 N28379 N28380 10
D28380 N28380 0 diode
R28381 N28380 N28381 10
D28381 N28381 0 diode
R28382 N28381 N28382 10
D28382 N28382 0 diode
R28383 N28382 N28383 10
D28383 N28383 0 diode
R28384 N28383 N28384 10
D28384 N28384 0 diode
R28385 N28384 N28385 10
D28385 N28385 0 diode
R28386 N28385 N28386 10
D28386 N28386 0 diode
R28387 N28386 N28387 10
D28387 N28387 0 diode
R28388 N28387 N28388 10
D28388 N28388 0 diode
R28389 N28388 N28389 10
D28389 N28389 0 diode
R28390 N28389 N28390 10
D28390 N28390 0 diode
R28391 N28390 N28391 10
D28391 N28391 0 diode
R28392 N28391 N28392 10
D28392 N28392 0 diode
R28393 N28392 N28393 10
D28393 N28393 0 diode
R28394 N28393 N28394 10
D28394 N28394 0 diode
R28395 N28394 N28395 10
D28395 N28395 0 diode
R28396 N28395 N28396 10
D28396 N28396 0 diode
R28397 N28396 N28397 10
D28397 N28397 0 diode
R28398 N28397 N28398 10
D28398 N28398 0 diode
R28399 N28398 N28399 10
D28399 N28399 0 diode
R28400 N28399 N28400 10
D28400 N28400 0 diode
R28401 N28400 N28401 10
D28401 N28401 0 diode
R28402 N28401 N28402 10
D28402 N28402 0 diode
R28403 N28402 N28403 10
D28403 N28403 0 diode
R28404 N28403 N28404 10
D28404 N28404 0 diode
R28405 N28404 N28405 10
D28405 N28405 0 diode
R28406 N28405 N28406 10
D28406 N28406 0 diode
R28407 N28406 N28407 10
D28407 N28407 0 diode
R28408 N28407 N28408 10
D28408 N28408 0 diode
R28409 N28408 N28409 10
D28409 N28409 0 diode
R28410 N28409 N28410 10
D28410 N28410 0 diode
R28411 N28410 N28411 10
D28411 N28411 0 diode
R28412 N28411 N28412 10
D28412 N28412 0 diode
R28413 N28412 N28413 10
D28413 N28413 0 diode
R28414 N28413 N28414 10
D28414 N28414 0 diode
R28415 N28414 N28415 10
D28415 N28415 0 diode
R28416 N28415 N28416 10
D28416 N28416 0 diode
R28417 N28416 N28417 10
D28417 N28417 0 diode
R28418 N28417 N28418 10
D28418 N28418 0 diode
R28419 N28418 N28419 10
D28419 N28419 0 diode
R28420 N28419 N28420 10
D28420 N28420 0 diode
R28421 N28420 N28421 10
D28421 N28421 0 diode
R28422 N28421 N28422 10
D28422 N28422 0 diode
R28423 N28422 N28423 10
D28423 N28423 0 diode
R28424 N28423 N28424 10
D28424 N28424 0 diode
R28425 N28424 N28425 10
D28425 N28425 0 diode
R28426 N28425 N28426 10
D28426 N28426 0 diode
R28427 N28426 N28427 10
D28427 N28427 0 diode
R28428 N28427 N28428 10
D28428 N28428 0 diode
R28429 N28428 N28429 10
D28429 N28429 0 diode
R28430 N28429 N28430 10
D28430 N28430 0 diode
R28431 N28430 N28431 10
D28431 N28431 0 diode
R28432 N28431 N28432 10
D28432 N28432 0 diode
R28433 N28432 N28433 10
D28433 N28433 0 diode
R28434 N28433 N28434 10
D28434 N28434 0 diode
R28435 N28434 N28435 10
D28435 N28435 0 diode
R28436 N28435 N28436 10
D28436 N28436 0 diode
R28437 N28436 N28437 10
D28437 N28437 0 diode
R28438 N28437 N28438 10
D28438 N28438 0 diode
R28439 N28438 N28439 10
D28439 N28439 0 diode
R28440 N28439 N28440 10
D28440 N28440 0 diode
R28441 N28440 N28441 10
D28441 N28441 0 diode
R28442 N28441 N28442 10
D28442 N28442 0 diode
R28443 N28442 N28443 10
D28443 N28443 0 diode
R28444 N28443 N28444 10
D28444 N28444 0 diode
R28445 N28444 N28445 10
D28445 N28445 0 diode
R28446 N28445 N28446 10
D28446 N28446 0 diode
R28447 N28446 N28447 10
D28447 N28447 0 diode
R28448 N28447 N28448 10
D28448 N28448 0 diode
R28449 N28448 N28449 10
D28449 N28449 0 diode
R28450 N28449 N28450 10
D28450 N28450 0 diode
R28451 N28450 N28451 10
D28451 N28451 0 diode
R28452 N28451 N28452 10
D28452 N28452 0 diode
R28453 N28452 N28453 10
D28453 N28453 0 diode
R28454 N28453 N28454 10
D28454 N28454 0 diode
R28455 N28454 N28455 10
D28455 N28455 0 diode
R28456 N28455 N28456 10
D28456 N28456 0 diode
R28457 N28456 N28457 10
D28457 N28457 0 diode
R28458 N28457 N28458 10
D28458 N28458 0 diode
R28459 N28458 N28459 10
D28459 N28459 0 diode
R28460 N28459 N28460 10
D28460 N28460 0 diode
R28461 N28460 N28461 10
D28461 N28461 0 diode
R28462 N28461 N28462 10
D28462 N28462 0 diode
R28463 N28462 N28463 10
D28463 N28463 0 diode
R28464 N28463 N28464 10
D28464 N28464 0 diode
R28465 N28464 N28465 10
D28465 N28465 0 diode
R28466 N28465 N28466 10
D28466 N28466 0 diode
R28467 N28466 N28467 10
D28467 N28467 0 diode
R28468 N28467 N28468 10
D28468 N28468 0 diode
R28469 N28468 N28469 10
D28469 N28469 0 diode
R28470 N28469 N28470 10
D28470 N28470 0 diode
R28471 N28470 N28471 10
D28471 N28471 0 diode
R28472 N28471 N28472 10
D28472 N28472 0 diode
R28473 N28472 N28473 10
D28473 N28473 0 diode
R28474 N28473 N28474 10
D28474 N28474 0 diode
R28475 N28474 N28475 10
D28475 N28475 0 diode
R28476 N28475 N28476 10
D28476 N28476 0 diode
R28477 N28476 N28477 10
D28477 N28477 0 diode
R28478 N28477 N28478 10
D28478 N28478 0 diode
R28479 N28478 N28479 10
D28479 N28479 0 diode
R28480 N28479 N28480 10
D28480 N28480 0 diode
R28481 N28480 N28481 10
D28481 N28481 0 diode
R28482 N28481 N28482 10
D28482 N28482 0 diode
R28483 N28482 N28483 10
D28483 N28483 0 diode
R28484 N28483 N28484 10
D28484 N28484 0 diode
R28485 N28484 N28485 10
D28485 N28485 0 diode
R28486 N28485 N28486 10
D28486 N28486 0 diode
R28487 N28486 N28487 10
D28487 N28487 0 diode
R28488 N28487 N28488 10
D28488 N28488 0 diode
R28489 N28488 N28489 10
D28489 N28489 0 diode
R28490 N28489 N28490 10
D28490 N28490 0 diode
R28491 N28490 N28491 10
D28491 N28491 0 diode
R28492 N28491 N28492 10
D28492 N28492 0 diode
R28493 N28492 N28493 10
D28493 N28493 0 diode
R28494 N28493 N28494 10
D28494 N28494 0 diode
R28495 N28494 N28495 10
D28495 N28495 0 diode
R28496 N28495 N28496 10
D28496 N28496 0 diode
R28497 N28496 N28497 10
D28497 N28497 0 diode
R28498 N28497 N28498 10
D28498 N28498 0 diode
R28499 N28498 N28499 10
D28499 N28499 0 diode
R28500 N28499 N28500 10
D28500 N28500 0 diode
R28501 N28500 N28501 10
D28501 N28501 0 diode
R28502 N28501 N28502 10
D28502 N28502 0 diode
R28503 N28502 N28503 10
D28503 N28503 0 diode
R28504 N28503 N28504 10
D28504 N28504 0 diode
R28505 N28504 N28505 10
D28505 N28505 0 diode
R28506 N28505 N28506 10
D28506 N28506 0 diode
R28507 N28506 N28507 10
D28507 N28507 0 diode
R28508 N28507 N28508 10
D28508 N28508 0 diode
R28509 N28508 N28509 10
D28509 N28509 0 diode
R28510 N28509 N28510 10
D28510 N28510 0 diode
R28511 N28510 N28511 10
D28511 N28511 0 diode
R28512 N28511 N28512 10
D28512 N28512 0 diode
R28513 N28512 N28513 10
D28513 N28513 0 diode
R28514 N28513 N28514 10
D28514 N28514 0 diode
R28515 N28514 N28515 10
D28515 N28515 0 diode
R28516 N28515 N28516 10
D28516 N28516 0 diode
R28517 N28516 N28517 10
D28517 N28517 0 diode
R28518 N28517 N28518 10
D28518 N28518 0 diode
R28519 N28518 N28519 10
D28519 N28519 0 diode
R28520 N28519 N28520 10
D28520 N28520 0 diode
R28521 N28520 N28521 10
D28521 N28521 0 diode
R28522 N28521 N28522 10
D28522 N28522 0 diode
R28523 N28522 N28523 10
D28523 N28523 0 diode
R28524 N28523 N28524 10
D28524 N28524 0 diode
R28525 N28524 N28525 10
D28525 N28525 0 diode
R28526 N28525 N28526 10
D28526 N28526 0 diode
R28527 N28526 N28527 10
D28527 N28527 0 diode
R28528 N28527 N28528 10
D28528 N28528 0 diode
R28529 N28528 N28529 10
D28529 N28529 0 diode
R28530 N28529 N28530 10
D28530 N28530 0 diode
R28531 N28530 N28531 10
D28531 N28531 0 diode
R28532 N28531 N28532 10
D28532 N28532 0 diode
R28533 N28532 N28533 10
D28533 N28533 0 diode
R28534 N28533 N28534 10
D28534 N28534 0 diode
R28535 N28534 N28535 10
D28535 N28535 0 diode
R28536 N28535 N28536 10
D28536 N28536 0 diode
R28537 N28536 N28537 10
D28537 N28537 0 diode
R28538 N28537 N28538 10
D28538 N28538 0 diode
R28539 N28538 N28539 10
D28539 N28539 0 diode
R28540 N28539 N28540 10
D28540 N28540 0 diode
R28541 N28540 N28541 10
D28541 N28541 0 diode
R28542 N28541 N28542 10
D28542 N28542 0 diode
R28543 N28542 N28543 10
D28543 N28543 0 diode
R28544 N28543 N28544 10
D28544 N28544 0 diode
R28545 N28544 N28545 10
D28545 N28545 0 diode
R28546 N28545 N28546 10
D28546 N28546 0 diode
R28547 N28546 N28547 10
D28547 N28547 0 diode
R28548 N28547 N28548 10
D28548 N28548 0 diode
R28549 N28548 N28549 10
D28549 N28549 0 diode
R28550 N28549 N28550 10
D28550 N28550 0 diode
R28551 N28550 N28551 10
D28551 N28551 0 diode
R28552 N28551 N28552 10
D28552 N28552 0 diode
R28553 N28552 N28553 10
D28553 N28553 0 diode
R28554 N28553 N28554 10
D28554 N28554 0 diode
R28555 N28554 N28555 10
D28555 N28555 0 diode
R28556 N28555 N28556 10
D28556 N28556 0 diode
R28557 N28556 N28557 10
D28557 N28557 0 diode
R28558 N28557 N28558 10
D28558 N28558 0 diode
R28559 N28558 N28559 10
D28559 N28559 0 diode
R28560 N28559 N28560 10
D28560 N28560 0 diode
R28561 N28560 N28561 10
D28561 N28561 0 diode
R28562 N28561 N28562 10
D28562 N28562 0 diode
R28563 N28562 N28563 10
D28563 N28563 0 diode
R28564 N28563 N28564 10
D28564 N28564 0 diode
R28565 N28564 N28565 10
D28565 N28565 0 diode
R28566 N28565 N28566 10
D28566 N28566 0 diode
R28567 N28566 N28567 10
D28567 N28567 0 diode
R28568 N28567 N28568 10
D28568 N28568 0 diode
R28569 N28568 N28569 10
D28569 N28569 0 diode
R28570 N28569 N28570 10
D28570 N28570 0 diode
R28571 N28570 N28571 10
D28571 N28571 0 diode
R28572 N28571 N28572 10
D28572 N28572 0 diode
R28573 N28572 N28573 10
D28573 N28573 0 diode
R28574 N28573 N28574 10
D28574 N28574 0 diode
R28575 N28574 N28575 10
D28575 N28575 0 diode
R28576 N28575 N28576 10
D28576 N28576 0 diode
R28577 N28576 N28577 10
D28577 N28577 0 diode
R28578 N28577 N28578 10
D28578 N28578 0 diode
R28579 N28578 N28579 10
D28579 N28579 0 diode
R28580 N28579 N28580 10
D28580 N28580 0 diode
R28581 N28580 N28581 10
D28581 N28581 0 diode
R28582 N28581 N28582 10
D28582 N28582 0 diode
R28583 N28582 N28583 10
D28583 N28583 0 diode
R28584 N28583 N28584 10
D28584 N28584 0 diode
R28585 N28584 N28585 10
D28585 N28585 0 diode
R28586 N28585 N28586 10
D28586 N28586 0 diode
R28587 N28586 N28587 10
D28587 N28587 0 diode
R28588 N28587 N28588 10
D28588 N28588 0 diode
R28589 N28588 N28589 10
D28589 N28589 0 diode
R28590 N28589 N28590 10
D28590 N28590 0 diode
R28591 N28590 N28591 10
D28591 N28591 0 diode
R28592 N28591 N28592 10
D28592 N28592 0 diode
R28593 N28592 N28593 10
D28593 N28593 0 diode
R28594 N28593 N28594 10
D28594 N28594 0 diode
R28595 N28594 N28595 10
D28595 N28595 0 diode
R28596 N28595 N28596 10
D28596 N28596 0 diode
R28597 N28596 N28597 10
D28597 N28597 0 diode
R28598 N28597 N28598 10
D28598 N28598 0 diode
R28599 N28598 N28599 10
D28599 N28599 0 diode
R28600 N28599 N28600 10
D28600 N28600 0 diode
R28601 N28600 N28601 10
D28601 N28601 0 diode
R28602 N28601 N28602 10
D28602 N28602 0 diode
R28603 N28602 N28603 10
D28603 N28603 0 diode
R28604 N28603 N28604 10
D28604 N28604 0 diode
R28605 N28604 N28605 10
D28605 N28605 0 diode
R28606 N28605 N28606 10
D28606 N28606 0 diode
R28607 N28606 N28607 10
D28607 N28607 0 diode
R28608 N28607 N28608 10
D28608 N28608 0 diode
R28609 N28608 N28609 10
D28609 N28609 0 diode
R28610 N28609 N28610 10
D28610 N28610 0 diode
R28611 N28610 N28611 10
D28611 N28611 0 diode
R28612 N28611 N28612 10
D28612 N28612 0 diode
R28613 N28612 N28613 10
D28613 N28613 0 diode
R28614 N28613 N28614 10
D28614 N28614 0 diode
R28615 N28614 N28615 10
D28615 N28615 0 diode
R28616 N28615 N28616 10
D28616 N28616 0 diode
R28617 N28616 N28617 10
D28617 N28617 0 diode
R28618 N28617 N28618 10
D28618 N28618 0 diode
R28619 N28618 N28619 10
D28619 N28619 0 diode
R28620 N28619 N28620 10
D28620 N28620 0 diode
R28621 N28620 N28621 10
D28621 N28621 0 diode
R28622 N28621 N28622 10
D28622 N28622 0 diode
R28623 N28622 N28623 10
D28623 N28623 0 diode
R28624 N28623 N28624 10
D28624 N28624 0 diode
R28625 N28624 N28625 10
D28625 N28625 0 diode
R28626 N28625 N28626 10
D28626 N28626 0 diode
R28627 N28626 N28627 10
D28627 N28627 0 diode
R28628 N28627 N28628 10
D28628 N28628 0 diode
R28629 N28628 N28629 10
D28629 N28629 0 diode
R28630 N28629 N28630 10
D28630 N28630 0 diode
R28631 N28630 N28631 10
D28631 N28631 0 diode
R28632 N28631 N28632 10
D28632 N28632 0 diode
R28633 N28632 N28633 10
D28633 N28633 0 diode
R28634 N28633 N28634 10
D28634 N28634 0 diode
R28635 N28634 N28635 10
D28635 N28635 0 diode
R28636 N28635 N28636 10
D28636 N28636 0 diode
R28637 N28636 N28637 10
D28637 N28637 0 diode
R28638 N28637 N28638 10
D28638 N28638 0 diode
R28639 N28638 N28639 10
D28639 N28639 0 diode
R28640 N28639 N28640 10
D28640 N28640 0 diode
R28641 N28640 N28641 10
D28641 N28641 0 diode
R28642 N28641 N28642 10
D28642 N28642 0 diode
R28643 N28642 N28643 10
D28643 N28643 0 diode
R28644 N28643 N28644 10
D28644 N28644 0 diode
R28645 N28644 N28645 10
D28645 N28645 0 diode
R28646 N28645 N28646 10
D28646 N28646 0 diode
R28647 N28646 N28647 10
D28647 N28647 0 diode
R28648 N28647 N28648 10
D28648 N28648 0 diode
R28649 N28648 N28649 10
D28649 N28649 0 diode
R28650 N28649 N28650 10
D28650 N28650 0 diode
R28651 N28650 N28651 10
D28651 N28651 0 diode
R28652 N28651 N28652 10
D28652 N28652 0 diode
R28653 N28652 N28653 10
D28653 N28653 0 diode
R28654 N28653 N28654 10
D28654 N28654 0 diode
R28655 N28654 N28655 10
D28655 N28655 0 diode
R28656 N28655 N28656 10
D28656 N28656 0 diode
R28657 N28656 N28657 10
D28657 N28657 0 diode
R28658 N28657 N28658 10
D28658 N28658 0 diode
R28659 N28658 N28659 10
D28659 N28659 0 diode
R28660 N28659 N28660 10
D28660 N28660 0 diode
R28661 N28660 N28661 10
D28661 N28661 0 diode
R28662 N28661 N28662 10
D28662 N28662 0 diode
R28663 N28662 N28663 10
D28663 N28663 0 diode
R28664 N28663 N28664 10
D28664 N28664 0 diode
R28665 N28664 N28665 10
D28665 N28665 0 diode
R28666 N28665 N28666 10
D28666 N28666 0 diode
R28667 N28666 N28667 10
D28667 N28667 0 diode
R28668 N28667 N28668 10
D28668 N28668 0 diode
R28669 N28668 N28669 10
D28669 N28669 0 diode
R28670 N28669 N28670 10
D28670 N28670 0 diode
R28671 N28670 N28671 10
D28671 N28671 0 diode
R28672 N28671 N28672 10
D28672 N28672 0 diode
R28673 N28672 N28673 10
D28673 N28673 0 diode
R28674 N28673 N28674 10
D28674 N28674 0 diode
R28675 N28674 N28675 10
D28675 N28675 0 diode
R28676 N28675 N28676 10
D28676 N28676 0 diode
R28677 N28676 N28677 10
D28677 N28677 0 diode
R28678 N28677 N28678 10
D28678 N28678 0 diode
R28679 N28678 N28679 10
D28679 N28679 0 diode
R28680 N28679 N28680 10
D28680 N28680 0 diode
R28681 N28680 N28681 10
D28681 N28681 0 diode
R28682 N28681 N28682 10
D28682 N28682 0 diode
R28683 N28682 N28683 10
D28683 N28683 0 diode
R28684 N28683 N28684 10
D28684 N28684 0 diode
R28685 N28684 N28685 10
D28685 N28685 0 diode
R28686 N28685 N28686 10
D28686 N28686 0 diode
R28687 N28686 N28687 10
D28687 N28687 0 diode
R28688 N28687 N28688 10
D28688 N28688 0 diode
R28689 N28688 N28689 10
D28689 N28689 0 diode
R28690 N28689 N28690 10
D28690 N28690 0 diode
R28691 N28690 N28691 10
D28691 N28691 0 diode
R28692 N28691 N28692 10
D28692 N28692 0 diode
R28693 N28692 N28693 10
D28693 N28693 0 diode
R28694 N28693 N28694 10
D28694 N28694 0 diode
R28695 N28694 N28695 10
D28695 N28695 0 diode
R28696 N28695 N28696 10
D28696 N28696 0 diode
R28697 N28696 N28697 10
D28697 N28697 0 diode
R28698 N28697 N28698 10
D28698 N28698 0 diode
R28699 N28698 N28699 10
D28699 N28699 0 diode
R28700 N28699 N28700 10
D28700 N28700 0 diode
R28701 N28700 N28701 10
D28701 N28701 0 diode
R28702 N28701 N28702 10
D28702 N28702 0 diode
R28703 N28702 N28703 10
D28703 N28703 0 diode
R28704 N28703 N28704 10
D28704 N28704 0 diode
R28705 N28704 N28705 10
D28705 N28705 0 diode
R28706 N28705 N28706 10
D28706 N28706 0 diode
R28707 N28706 N28707 10
D28707 N28707 0 diode
R28708 N28707 N28708 10
D28708 N28708 0 diode
R28709 N28708 N28709 10
D28709 N28709 0 diode
R28710 N28709 N28710 10
D28710 N28710 0 diode
R28711 N28710 N28711 10
D28711 N28711 0 diode
R28712 N28711 N28712 10
D28712 N28712 0 diode
R28713 N28712 N28713 10
D28713 N28713 0 diode
R28714 N28713 N28714 10
D28714 N28714 0 diode
R28715 N28714 N28715 10
D28715 N28715 0 diode
R28716 N28715 N28716 10
D28716 N28716 0 diode
R28717 N28716 N28717 10
D28717 N28717 0 diode
R28718 N28717 N28718 10
D28718 N28718 0 diode
R28719 N28718 N28719 10
D28719 N28719 0 diode
R28720 N28719 N28720 10
D28720 N28720 0 diode
R28721 N28720 N28721 10
D28721 N28721 0 diode
R28722 N28721 N28722 10
D28722 N28722 0 diode
R28723 N28722 N28723 10
D28723 N28723 0 diode
R28724 N28723 N28724 10
D28724 N28724 0 diode
R28725 N28724 N28725 10
D28725 N28725 0 diode
R28726 N28725 N28726 10
D28726 N28726 0 diode
R28727 N28726 N28727 10
D28727 N28727 0 diode
R28728 N28727 N28728 10
D28728 N28728 0 diode
R28729 N28728 N28729 10
D28729 N28729 0 diode
R28730 N28729 N28730 10
D28730 N28730 0 diode
R28731 N28730 N28731 10
D28731 N28731 0 diode
R28732 N28731 N28732 10
D28732 N28732 0 diode
R28733 N28732 N28733 10
D28733 N28733 0 diode
R28734 N28733 N28734 10
D28734 N28734 0 diode
R28735 N28734 N28735 10
D28735 N28735 0 diode
R28736 N28735 N28736 10
D28736 N28736 0 diode
R28737 N28736 N28737 10
D28737 N28737 0 diode
R28738 N28737 N28738 10
D28738 N28738 0 diode
R28739 N28738 N28739 10
D28739 N28739 0 diode
R28740 N28739 N28740 10
D28740 N28740 0 diode
R28741 N28740 N28741 10
D28741 N28741 0 diode
R28742 N28741 N28742 10
D28742 N28742 0 diode
R28743 N28742 N28743 10
D28743 N28743 0 diode
R28744 N28743 N28744 10
D28744 N28744 0 diode
R28745 N28744 N28745 10
D28745 N28745 0 diode
R28746 N28745 N28746 10
D28746 N28746 0 diode
R28747 N28746 N28747 10
D28747 N28747 0 diode
R28748 N28747 N28748 10
D28748 N28748 0 diode
R28749 N28748 N28749 10
D28749 N28749 0 diode
R28750 N28749 N28750 10
D28750 N28750 0 diode
R28751 N28750 N28751 10
D28751 N28751 0 diode
R28752 N28751 N28752 10
D28752 N28752 0 diode
R28753 N28752 N28753 10
D28753 N28753 0 diode
R28754 N28753 N28754 10
D28754 N28754 0 diode
R28755 N28754 N28755 10
D28755 N28755 0 diode
R28756 N28755 N28756 10
D28756 N28756 0 diode
R28757 N28756 N28757 10
D28757 N28757 0 diode
R28758 N28757 N28758 10
D28758 N28758 0 diode
R28759 N28758 N28759 10
D28759 N28759 0 diode
R28760 N28759 N28760 10
D28760 N28760 0 diode
R28761 N28760 N28761 10
D28761 N28761 0 diode
R28762 N28761 N28762 10
D28762 N28762 0 diode
R28763 N28762 N28763 10
D28763 N28763 0 diode
R28764 N28763 N28764 10
D28764 N28764 0 diode
R28765 N28764 N28765 10
D28765 N28765 0 diode
R28766 N28765 N28766 10
D28766 N28766 0 diode
R28767 N28766 N28767 10
D28767 N28767 0 diode
R28768 N28767 N28768 10
D28768 N28768 0 diode
R28769 N28768 N28769 10
D28769 N28769 0 diode
R28770 N28769 N28770 10
D28770 N28770 0 diode
R28771 N28770 N28771 10
D28771 N28771 0 diode
R28772 N28771 N28772 10
D28772 N28772 0 diode
R28773 N28772 N28773 10
D28773 N28773 0 diode
R28774 N28773 N28774 10
D28774 N28774 0 diode
R28775 N28774 N28775 10
D28775 N28775 0 diode
R28776 N28775 N28776 10
D28776 N28776 0 diode
R28777 N28776 N28777 10
D28777 N28777 0 diode
R28778 N28777 N28778 10
D28778 N28778 0 diode
R28779 N28778 N28779 10
D28779 N28779 0 diode
R28780 N28779 N28780 10
D28780 N28780 0 diode
R28781 N28780 N28781 10
D28781 N28781 0 diode
R28782 N28781 N28782 10
D28782 N28782 0 diode
R28783 N28782 N28783 10
D28783 N28783 0 diode
R28784 N28783 N28784 10
D28784 N28784 0 diode
R28785 N28784 N28785 10
D28785 N28785 0 diode
R28786 N28785 N28786 10
D28786 N28786 0 diode
R28787 N28786 N28787 10
D28787 N28787 0 diode
R28788 N28787 N28788 10
D28788 N28788 0 diode
R28789 N28788 N28789 10
D28789 N28789 0 diode
R28790 N28789 N28790 10
D28790 N28790 0 diode
R28791 N28790 N28791 10
D28791 N28791 0 diode
R28792 N28791 N28792 10
D28792 N28792 0 diode
R28793 N28792 N28793 10
D28793 N28793 0 diode
R28794 N28793 N28794 10
D28794 N28794 0 diode
R28795 N28794 N28795 10
D28795 N28795 0 diode
R28796 N28795 N28796 10
D28796 N28796 0 diode
R28797 N28796 N28797 10
D28797 N28797 0 diode
R28798 N28797 N28798 10
D28798 N28798 0 diode
R28799 N28798 N28799 10
D28799 N28799 0 diode
R28800 N28799 N28800 10
D28800 N28800 0 diode
R28801 N28800 N28801 10
D28801 N28801 0 diode
R28802 N28801 N28802 10
D28802 N28802 0 diode
R28803 N28802 N28803 10
D28803 N28803 0 diode
R28804 N28803 N28804 10
D28804 N28804 0 diode
R28805 N28804 N28805 10
D28805 N28805 0 diode
R28806 N28805 N28806 10
D28806 N28806 0 diode
R28807 N28806 N28807 10
D28807 N28807 0 diode
R28808 N28807 N28808 10
D28808 N28808 0 diode
R28809 N28808 N28809 10
D28809 N28809 0 diode
R28810 N28809 N28810 10
D28810 N28810 0 diode
R28811 N28810 N28811 10
D28811 N28811 0 diode
R28812 N28811 N28812 10
D28812 N28812 0 diode
R28813 N28812 N28813 10
D28813 N28813 0 diode
R28814 N28813 N28814 10
D28814 N28814 0 diode
R28815 N28814 N28815 10
D28815 N28815 0 diode
R28816 N28815 N28816 10
D28816 N28816 0 diode
R28817 N28816 N28817 10
D28817 N28817 0 diode
R28818 N28817 N28818 10
D28818 N28818 0 diode
R28819 N28818 N28819 10
D28819 N28819 0 diode
R28820 N28819 N28820 10
D28820 N28820 0 diode
R28821 N28820 N28821 10
D28821 N28821 0 diode
R28822 N28821 N28822 10
D28822 N28822 0 diode
R28823 N28822 N28823 10
D28823 N28823 0 diode
R28824 N28823 N28824 10
D28824 N28824 0 diode
R28825 N28824 N28825 10
D28825 N28825 0 diode
R28826 N28825 N28826 10
D28826 N28826 0 diode
R28827 N28826 N28827 10
D28827 N28827 0 diode
R28828 N28827 N28828 10
D28828 N28828 0 diode
R28829 N28828 N28829 10
D28829 N28829 0 diode
R28830 N28829 N28830 10
D28830 N28830 0 diode
R28831 N28830 N28831 10
D28831 N28831 0 diode
R28832 N28831 N28832 10
D28832 N28832 0 diode
R28833 N28832 N28833 10
D28833 N28833 0 diode
R28834 N28833 N28834 10
D28834 N28834 0 diode
R28835 N28834 N28835 10
D28835 N28835 0 diode
R28836 N28835 N28836 10
D28836 N28836 0 diode
R28837 N28836 N28837 10
D28837 N28837 0 diode
R28838 N28837 N28838 10
D28838 N28838 0 diode
R28839 N28838 N28839 10
D28839 N28839 0 diode
R28840 N28839 N28840 10
D28840 N28840 0 diode
R28841 N28840 N28841 10
D28841 N28841 0 diode
R28842 N28841 N28842 10
D28842 N28842 0 diode
R28843 N28842 N28843 10
D28843 N28843 0 diode
R28844 N28843 N28844 10
D28844 N28844 0 diode
R28845 N28844 N28845 10
D28845 N28845 0 diode
R28846 N28845 N28846 10
D28846 N28846 0 diode
R28847 N28846 N28847 10
D28847 N28847 0 diode
R28848 N28847 N28848 10
D28848 N28848 0 diode
R28849 N28848 N28849 10
D28849 N28849 0 diode
R28850 N28849 N28850 10
D28850 N28850 0 diode
R28851 N28850 N28851 10
D28851 N28851 0 diode
R28852 N28851 N28852 10
D28852 N28852 0 diode
R28853 N28852 N28853 10
D28853 N28853 0 diode
R28854 N28853 N28854 10
D28854 N28854 0 diode
R28855 N28854 N28855 10
D28855 N28855 0 diode
R28856 N28855 N28856 10
D28856 N28856 0 diode
R28857 N28856 N28857 10
D28857 N28857 0 diode
R28858 N28857 N28858 10
D28858 N28858 0 diode
R28859 N28858 N28859 10
D28859 N28859 0 diode
R28860 N28859 N28860 10
D28860 N28860 0 diode
R28861 N28860 N28861 10
D28861 N28861 0 diode
R28862 N28861 N28862 10
D28862 N28862 0 diode
R28863 N28862 N28863 10
D28863 N28863 0 diode
R28864 N28863 N28864 10
D28864 N28864 0 diode
R28865 N28864 N28865 10
D28865 N28865 0 diode
R28866 N28865 N28866 10
D28866 N28866 0 diode
R28867 N28866 N28867 10
D28867 N28867 0 diode
R28868 N28867 N28868 10
D28868 N28868 0 diode
R28869 N28868 N28869 10
D28869 N28869 0 diode
R28870 N28869 N28870 10
D28870 N28870 0 diode
R28871 N28870 N28871 10
D28871 N28871 0 diode
R28872 N28871 N28872 10
D28872 N28872 0 diode
R28873 N28872 N28873 10
D28873 N28873 0 diode
R28874 N28873 N28874 10
D28874 N28874 0 diode
R28875 N28874 N28875 10
D28875 N28875 0 diode
R28876 N28875 N28876 10
D28876 N28876 0 diode
R28877 N28876 N28877 10
D28877 N28877 0 diode
R28878 N28877 N28878 10
D28878 N28878 0 diode
R28879 N28878 N28879 10
D28879 N28879 0 diode
R28880 N28879 N28880 10
D28880 N28880 0 diode
R28881 N28880 N28881 10
D28881 N28881 0 diode
R28882 N28881 N28882 10
D28882 N28882 0 diode
R28883 N28882 N28883 10
D28883 N28883 0 diode
R28884 N28883 N28884 10
D28884 N28884 0 diode
R28885 N28884 N28885 10
D28885 N28885 0 diode
R28886 N28885 N28886 10
D28886 N28886 0 diode
R28887 N28886 N28887 10
D28887 N28887 0 diode
R28888 N28887 N28888 10
D28888 N28888 0 diode
R28889 N28888 N28889 10
D28889 N28889 0 diode
R28890 N28889 N28890 10
D28890 N28890 0 diode
R28891 N28890 N28891 10
D28891 N28891 0 diode
R28892 N28891 N28892 10
D28892 N28892 0 diode
R28893 N28892 N28893 10
D28893 N28893 0 diode
R28894 N28893 N28894 10
D28894 N28894 0 diode
R28895 N28894 N28895 10
D28895 N28895 0 diode
R28896 N28895 N28896 10
D28896 N28896 0 diode
R28897 N28896 N28897 10
D28897 N28897 0 diode
R28898 N28897 N28898 10
D28898 N28898 0 diode
R28899 N28898 N28899 10
D28899 N28899 0 diode
R28900 N28899 N28900 10
D28900 N28900 0 diode
R28901 N28900 N28901 10
D28901 N28901 0 diode
R28902 N28901 N28902 10
D28902 N28902 0 diode
R28903 N28902 N28903 10
D28903 N28903 0 diode
R28904 N28903 N28904 10
D28904 N28904 0 diode
R28905 N28904 N28905 10
D28905 N28905 0 diode
R28906 N28905 N28906 10
D28906 N28906 0 diode
R28907 N28906 N28907 10
D28907 N28907 0 diode
R28908 N28907 N28908 10
D28908 N28908 0 diode
R28909 N28908 N28909 10
D28909 N28909 0 diode
R28910 N28909 N28910 10
D28910 N28910 0 diode
R28911 N28910 N28911 10
D28911 N28911 0 diode
R28912 N28911 N28912 10
D28912 N28912 0 diode
R28913 N28912 N28913 10
D28913 N28913 0 diode
R28914 N28913 N28914 10
D28914 N28914 0 diode
R28915 N28914 N28915 10
D28915 N28915 0 diode
R28916 N28915 N28916 10
D28916 N28916 0 diode
R28917 N28916 N28917 10
D28917 N28917 0 diode
R28918 N28917 N28918 10
D28918 N28918 0 diode
R28919 N28918 N28919 10
D28919 N28919 0 diode
R28920 N28919 N28920 10
D28920 N28920 0 diode
R28921 N28920 N28921 10
D28921 N28921 0 diode
R28922 N28921 N28922 10
D28922 N28922 0 diode
R28923 N28922 N28923 10
D28923 N28923 0 diode
R28924 N28923 N28924 10
D28924 N28924 0 diode
R28925 N28924 N28925 10
D28925 N28925 0 diode
R28926 N28925 N28926 10
D28926 N28926 0 diode
R28927 N28926 N28927 10
D28927 N28927 0 diode
R28928 N28927 N28928 10
D28928 N28928 0 diode
R28929 N28928 N28929 10
D28929 N28929 0 diode
R28930 N28929 N28930 10
D28930 N28930 0 diode
R28931 N28930 N28931 10
D28931 N28931 0 diode
R28932 N28931 N28932 10
D28932 N28932 0 diode
R28933 N28932 N28933 10
D28933 N28933 0 diode
R28934 N28933 N28934 10
D28934 N28934 0 diode
R28935 N28934 N28935 10
D28935 N28935 0 diode
R28936 N28935 N28936 10
D28936 N28936 0 diode
R28937 N28936 N28937 10
D28937 N28937 0 diode
R28938 N28937 N28938 10
D28938 N28938 0 diode
R28939 N28938 N28939 10
D28939 N28939 0 diode
R28940 N28939 N28940 10
D28940 N28940 0 diode
R28941 N28940 N28941 10
D28941 N28941 0 diode
R28942 N28941 N28942 10
D28942 N28942 0 diode
R28943 N28942 N28943 10
D28943 N28943 0 diode
R28944 N28943 N28944 10
D28944 N28944 0 diode
R28945 N28944 N28945 10
D28945 N28945 0 diode
R28946 N28945 N28946 10
D28946 N28946 0 diode
R28947 N28946 N28947 10
D28947 N28947 0 diode
R28948 N28947 N28948 10
D28948 N28948 0 diode
R28949 N28948 N28949 10
D28949 N28949 0 diode
R28950 N28949 N28950 10
D28950 N28950 0 diode
R28951 N28950 N28951 10
D28951 N28951 0 diode
R28952 N28951 N28952 10
D28952 N28952 0 diode
R28953 N28952 N28953 10
D28953 N28953 0 diode
R28954 N28953 N28954 10
D28954 N28954 0 diode
R28955 N28954 N28955 10
D28955 N28955 0 diode
R28956 N28955 N28956 10
D28956 N28956 0 diode
R28957 N28956 N28957 10
D28957 N28957 0 diode
R28958 N28957 N28958 10
D28958 N28958 0 diode
R28959 N28958 N28959 10
D28959 N28959 0 diode
R28960 N28959 N28960 10
D28960 N28960 0 diode
R28961 N28960 N28961 10
D28961 N28961 0 diode
R28962 N28961 N28962 10
D28962 N28962 0 diode
R28963 N28962 N28963 10
D28963 N28963 0 diode
R28964 N28963 N28964 10
D28964 N28964 0 diode
R28965 N28964 N28965 10
D28965 N28965 0 diode
R28966 N28965 N28966 10
D28966 N28966 0 diode
R28967 N28966 N28967 10
D28967 N28967 0 diode
R28968 N28967 N28968 10
D28968 N28968 0 diode
R28969 N28968 N28969 10
D28969 N28969 0 diode
R28970 N28969 N28970 10
D28970 N28970 0 diode
R28971 N28970 N28971 10
D28971 N28971 0 diode
R28972 N28971 N28972 10
D28972 N28972 0 diode
R28973 N28972 N28973 10
D28973 N28973 0 diode
R28974 N28973 N28974 10
D28974 N28974 0 diode
R28975 N28974 N28975 10
D28975 N28975 0 diode
R28976 N28975 N28976 10
D28976 N28976 0 diode
R28977 N28976 N28977 10
D28977 N28977 0 diode
R28978 N28977 N28978 10
D28978 N28978 0 diode
R28979 N28978 N28979 10
D28979 N28979 0 diode
R28980 N28979 N28980 10
D28980 N28980 0 diode
R28981 N28980 N28981 10
D28981 N28981 0 diode
R28982 N28981 N28982 10
D28982 N28982 0 diode
R28983 N28982 N28983 10
D28983 N28983 0 diode
R28984 N28983 N28984 10
D28984 N28984 0 diode
R28985 N28984 N28985 10
D28985 N28985 0 diode
R28986 N28985 N28986 10
D28986 N28986 0 diode
R28987 N28986 N28987 10
D28987 N28987 0 diode
R28988 N28987 N28988 10
D28988 N28988 0 diode
R28989 N28988 N28989 10
D28989 N28989 0 diode
R28990 N28989 N28990 10
D28990 N28990 0 diode
R28991 N28990 N28991 10
D28991 N28991 0 diode
R28992 N28991 N28992 10
D28992 N28992 0 diode
R28993 N28992 N28993 10
D28993 N28993 0 diode
R28994 N28993 N28994 10
D28994 N28994 0 diode
R28995 N28994 N28995 10
D28995 N28995 0 diode
R28996 N28995 N28996 10
D28996 N28996 0 diode
R28997 N28996 N28997 10
D28997 N28997 0 diode
R28998 N28997 N28998 10
D28998 N28998 0 diode
R28999 N28998 N28999 10
D28999 N28999 0 diode
R29000 N28999 N29000 10
D29000 N29000 0 diode
R29001 N29000 N29001 10
D29001 N29001 0 diode
R29002 N29001 N29002 10
D29002 N29002 0 diode
R29003 N29002 N29003 10
D29003 N29003 0 diode
R29004 N29003 N29004 10
D29004 N29004 0 diode
R29005 N29004 N29005 10
D29005 N29005 0 diode
R29006 N29005 N29006 10
D29006 N29006 0 diode
R29007 N29006 N29007 10
D29007 N29007 0 diode
R29008 N29007 N29008 10
D29008 N29008 0 diode
R29009 N29008 N29009 10
D29009 N29009 0 diode
R29010 N29009 N29010 10
D29010 N29010 0 diode
R29011 N29010 N29011 10
D29011 N29011 0 diode
R29012 N29011 N29012 10
D29012 N29012 0 diode
R29013 N29012 N29013 10
D29013 N29013 0 diode
R29014 N29013 N29014 10
D29014 N29014 0 diode
R29015 N29014 N29015 10
D29015 N29015 0 diode
R29016 N29015 N29016 10
D29016 N29016 0 diode
R29017 N29016 N29017 10
D29017 N29017 0 diode
R29018 N29017 N29018 10
D29018 N29018 0 diode
R29019 N29018 N29019 10
D29019 N29019 0 diode
R29020 N29019 N29020 10
D29020 N29020 0 diode
R29021 N29020 N29021 10
D29021 N29021 0 diode
R29022 N29021 N29022 10
D29022 N29022 0 diode
R29023 N29022 N29023 10
D29023 N29023 0 diode
R29024 N29023 N29024 10
D29024 N29024 0 diode
R29025 N29024 N29025 10
D29025 N29025 0 diode
R29026 N29025 N29026 10
D29026 N29026 0 diode
R29027 N29026 N29027 10
D29027 N29027 0 diode
R29028 N29027 N29028 10
D29028 N29028 0 diode
R29029 N29028 N29029 10
D29029 N29029 0 diode
R29030 N29029 N29030 10
D29030 N29030 0 diode
R29031 N29030 N29031 10
D29031 N29031 0 diode
R29032 N29031 N29032 10
D29032 N29032 0 diode
R29033 N29032 N29033 10
D29033 N29033 0 diode
R29034 N29033 N29034 10
D29034 N29034 0 diode
R29035 N29034 N29035 10
D29035 N29035 0 diode
R29036 N29035 N29036 10
D29036 N29036 0 diode
R29037 N29036 N29037 10
D29037 N29037 0 diode
R29038 N29037 N29038 10
D29038 N29038 0 diode
R29039 N29038 N29039 10
D29039 N29039 0 diode
R29040 N29039 N29040 10
D29040 N29040 0 diode
R29041 N29040 N29041 10
D29041 N29041 0 diode
R29042 N29041 N29042 10
D29042 N29042 0 diode
R29043 N29042 N29043 10
D29043 N29043 0 diode
R29044 N29043 N29044 10
D29044 N29044 0 diode
R29045 N29044 N29045 10
D29045 N29045 0 diode
R29046 N29045 N29046 10
D29046 N29046 0 diode
R29047 N29046 N29047 10
D29047 N29047 0 diode
R29048 N29047 N29048 10
D29048 N29048 0 diode
R29049 N29048 N29049 10
D29049 N29049 0 diode
R29050 N29049 N29050 10
D29050 N29050 0 diode
R29051 N29050 N29051 10
D29051 N29051 0 diode
R29052 N29051 N29052 10
D29052 N29052 0 diode
R29053 N29052 N29053 10
D29053 N29053 0 diode
R29054 N29053 N29054 10
D29054 N29054 0 diode
R29055 N29054 N29055 10
D29055 N29055 0 diode
R29056 N29055 N29056 10
D29056 N29056 0 diode
R29057 N29056 N29057 10
D29057 N29057 0 diode
R29058 N29057 N29058 10
D29058 N29058 0 diode
R29059 N29058 N29059 10
D29059 N29059 0 diode
R29060 N29059 N29060 10
D29060 N29060 0 diode
R29061 N29060 N29061 10
D29061 N29061 0 diode
R29062 N29061 N29062 10
D29062 N29062 0 diode
R29063 N29062 N29063 10
D29063 N29063 0 diode
R29064 N29063 N29064 10
D29064 N29064 0 diode
R29065 N29064 N29065 10
D29065 N29065 0 diode
R29066 N29065 N29066 10
D29066 N29066 0 diode
R29067 N29066 N29067 10
D29067 N29067 0 diode
R29068 N29067 N29068 10
D29068 N29068 0 diode
R29069 N29068 N29069 10
D29069 N29069 0 diode
R29070 N29069 N29070 10
D29070 N29070 0 diode
R29071 N29070 N29071 10
D29071 N29071 0 diode
R29072 N29071 N29072 10
D29072 N29072 0 diode
R29073 N29072 N29073 10
D29073 N29073 0 diode
R29074 N29073 N29074 10
D29074 N29074 0 diode
R29075 N29074 N29075 10
D29075 N29075 0 diode
R29076 N29075 N29076 10
D29076 N29076 0 diode
R29077 N29076 N29077 10
D29077 N29077 0 diode
R29078 N29077 N29078 10
D29078 N29078 0 diode
R29079 N29078 N29079 10
D29079 N29079 0 diode
R29080 N29079 N29080 10
D29080 N29080 0 diode
R29081 N29080 N29081 10
D29081 N29081 0 diode
R29082 N29081 N29082 10
D29082 N29082 0 diode
R29083 N29082 N29083 10
D29083 N29083 0 diode
R29084 N29083 N29084 10
D29084 N29084 0 diode
R29085 N29084 N29085 10
D29085 N29085 0 diode
R29086 N29085 N29086 10
D29086 N29086 0 diode
R29087 N29086 N29087 10
D29087 N29087 0 diode
R29088 N29087 N29088 10
D29088 N29088 0 diode
R29089 N29088 N29089 10
D29089 N29089 0 diode
R29090 N29089 N29090 10
D29090 N29090 0 diode
R29091 N29090 N29091 10
D29091 N29091 0 diode
R29092 N29091 N29092 10
D29092 N29092 0 diode
R29093 N29092 N29093 10
D29093 N29093 0 diode
R29094 N29093 N29094 10
D29094 N29094 0 diode
R29095 N29094 N29095 10
D29095 N29095 0 diode
R29096 N29095 N29096 10
D29096 N29096 0 diode
R29097 N29096 N29097 10
D29097 N29097 0 diode
R29098 N29097 N29098 10
D29098 N29098 0 diode
R29099 N29098 N29099 10
D29099 N29099 0 diode
R29100 N29099 N29100 10
D29100 N29100 0 diode
R29101 N29100 N29101 10
D29101 N29101 0 diode
R29102 N29101 N29102 10
D29102 N29102 0 diode
R29103 N29102 N29103 10
D29103 N29103 0 diode
R29104 N29103 N29104 10
D29104 N29104 0 diode
R29105 N29104 N29105 10
D29105 N29105 0 diode
R29106 N29105 N29106 10
D29106 N29106 0 diode
R29107 N29106 N29107 10
D29107 N29107 0 diode
R29108 N29107 N29108 10
D29108 N29108 0 diode
R29109 N29108 N29109 10
D29109 N29109 0 diode
R29110 N29109 N29110 10
D29110 N29110 0 diode
R29111 N29110 N29111 10
D29111 N29111 0 diode
R29112 N29111 N29112 10
D29112 N29112 0 diode
R29113 N29112 N29113 10
D29113 N29113 0 diode
R29114 N29113 N29114 10
D29114 N29114 0 diode
R29115 N29114 N29115 10
D29115 N29115 0 diode
R29116 N29115 N29116 10
D29116 N29116 0 diode
R29117 N29116 N29117 10
D29117 N29117 0 diode
R29118 N29117 N29118 10
D29118 N29118 0 diode
R29119 N29118 N29119 10
D29119 N29119 0 diode
R29120 N29119 N29120 10
D29120 N29120 0 diode
R29121 N29120 N29121 10
D29121 N29121 0 diode
R29122 N29121 N29122 10
D29122 N29122 0 diode
R29123 N29122 N29123 10
D29123 N29123 0 diode
R29124 N29123 N29124 10
D29124 N29124 0 diode
R29125 N29124 N29125 10
D29125 N29125 0 diode
R29126 N29125 N29126 10
D29126 N29126 0 diode
R29127 N29126 N29127 10
D29127 N29127 0 diode
R29128 N29127 N29128 10
D29128 N29128 0 diode
R29129 N29128 N29129 10
D29129 N29129 0 diode
R29130 N29129 N29130 10
D29130 N29130 0 diode
R29131 N29130 N29131 10
D29131 N29131 0 diode
R29132 N29131 N29132 10
D29132 N29132 0 diode
R29133 N29132 N29133 10
D29133 N29133 0 diode
R29134 N29133 N29134 10
D29134 N29134 0 diode
R29135 N29134 N29135 10
D29135 N29135 0 diode
R29136 N29135 N29136 10
D29136 N29136 0 diode
R29137 N29136 N29137 10
D29137 N29137 0 diode
R29138 N29137 N29138 10
D29138 N29138 0 diode
R29139 N29138 N29139 10
D29139 N29139 0 diode
R29140 N29139 N29140 10
D29140 N29140 0 diode
R29141 N29140 N29141 10
D29141 N29141 0 diode
R29142 N29141 N29142 10
D29142 N29142 0 diode
R29143 N29142 N29143 10
D29143 N29143 0 diode
R29144 N29143 N29144 10
D29144 N29144 0 diode
R29145 N29144 N29145 10
D29145 N29145 0 diode
R29146 N29145 N29146 10
D29146 N29146 0 diode
R29147 N29146 N29147 10
D29147 N29147 0 diode
R29148 N29147 N29148 10
D29148 N29148 0 diode
R29149 N29148 N29149 10
D29149 N29149 0 diode
R29150 N29149 N29150 10
D29150 N29150 0 diode
R29151 N29150 N29151 10
D29151 N29151 0 diode
R29152 N29151 N29152 10
D29152 N29152 0 diode
R29153 N29152 N29153 10
D29153 N29153 0 diode
R29154 N29153 N29154 10
D29154 N29154 0 diode
R29155 N29154 N29155 10
D29155 N29155 0 diode
R29156 N29155 N29156 10
D29156 N29156 0 diode
R29157 N29156 N29157 10
D29157 N29157 0 diode
R29158 N29157 N29158 10
D29158 N29158 0 diode
R29159 N29158 N29159 10
D29159 N29159 0 diode
R29160 N29159 N29160 10
D29160 N29160 0 diode
R29161 N29160 N29161 10
D29161 N29161 0 diode
R29162 N29161 N29162 10
D29162 N29162 0 diode
R29163 N29162 N29163 10
D29163 N29163 0 diode
R29164 N29163 N29164 10
D29164 N29164 0 diode
R29165 N29164 N29165 10
D29165 N29165 0 diode
R29166 N29165 N29166 10
D29166 N29166 0 diode
R29167 N29166 N29167 10
D29167 N29167 0 diode
R29168 N29167 N29168 10
D29168 N29168 0 diode
R29169 N29168 N29169 10
D29169 N29169 0 diode
R29170 N29169 N29170 10
D29170 N29170 0 diode
R29171 N29170 N29171 10
D29171 N29171 0 diode
R29172 N29171 N29172 10
D29172 N29172 0 diode
R29173 N29172 N29173 10
D29173 N29173 0 diode
R29174 N29173 N29174 10
D29174 N29174 0 diode
R29175 N29174 N29175 10
D29175 N29175 0 diode
R29176 N29175 N29176 10
D29176 N29176 0 diode
R29177 N29176 N29177 10
D29177 N29177 0 diode
R29178 N29177 N29178 10
D29178 N29178 0 diode
R29179 N29178 N29179 10
D29179 N29179 0 diode
R29180 N29179 N29180 10
D29180 N29180 0 diode
R29181 N29180 N29181 10
D29181 N29181 0 diode
R29182 N29181 N29182 10
D29182 N29182 0 diode
R29183 N29182 N29183 10
D29183 N29183 0 diode
R29184 N29183 N29184 10
D29184 N29184 0 diode
R29185 N29184 N29185 10
D29185 N29185 0 diode
R29186 N29185 N29186 10
D29186 N29186 0 diode
R29187 N29186 N29187 10
D29187 N29187 0 diode
R29188 N29187 N29188 10
D29188 N29188 0 diode
R29189 N29188 N29189 10
D29189 N29189 0 diode
R29190 N29189 N29190 10
D29190 N29190 0 diode
R29191 N29190 N29191 10
D29191 N29191 0 diode
R29192 N29191 N29192 10
D29192 N29192 0 diode
R29193 N29192 N29193 10
D29193 N29193 0 diode
R29194 N29193 N29194 10
D29194 N29194 0 diode
R29195 N29194 N29195 10
D29195 N29195 0 diode
R29196 N29195 N29196 10
D29196 N29196 0 diode
R29197 N29196 N29197 10
D29197 N29197 0 diode
R29198 N29197 N29198 10
D29198 N29198 0 diode
R29199 N29198 N29199 10
D29199 N29199 0 diode
R29200 N29199 N29200 10
D29200 N29200 0 diode
R29201 N29200 N29201 10
D29201 N29201 0 diode
R29202 N29201 N29202 10
D29202 N29202 0 diode
R29203 N29202 N29203 10
D29203 N29203 0 diode
R29204 N29203 N29204 10
D29204 N29204 0 diode
R29205 N29204 N29205 10
D29205 N29205 0 diode
R29206 N29205 N29206 10
D29206 N29206 0 diode
R29207 N29206 N29207 10
D29207 N29207 0 diode
R29208 N29207 N29208 10
D29208 N29208 0 diode
R29209 N29208 N29209 10
D29209 N29209 0 diode
R29210 N29209 N29210 10
D29210 N29210 0 diode
R29211 N29210 N29211 10
D29211 N29211 0 diode
R29212 N29211 N29212 10
D29212 N29212 0 diode
R29213 N29212 N29213 10
D29213 N29213 0 diode
R29214 N29213 N29214 10
D29214 N29214 0 diode
R29215 N29214 N29215 10
D29215 N29215 0 diode
R29216 N29215 N29216 10
D29216 N29216 0 diode
R29217 N29216 N29217 10
D29217 N29217 0 diode
R29218 N29217 N29218 10
D29218 N29218 0 diode
R29219 N29218 N29219 10
D29219 N29219 0 diode
R29220 N29219 N29220 10
D29220 N29220 0 diode
R29221 N29220 N29221 10
D29221 N29221 0 diode
R29222 N29221 N29222 10
D29222 N29222 0 diode
R29223 N29222 N29223 10
D29223 N29223 0 diode
R29224 N29223 N29224 10
D29224 N29224 0 diode
R29225 N29224 N29225 10
D29225 N29225 0 diode
R29226 N29225 N29226 10
D29226 N29226 0 diode
R29227 N29226 N29227 10
D29227 N29227 0 diode
R29228 N29227 N29228 10
D29228 N29228 0 diode
R29229 N29228 N29229 10
D29229 N29229 0 diode
R29230 N29229 N29230 10
D29230 N29230 0 diode
R29231 N29230 N29231 10
D29231 N29231 0 diode
R29232 N29231 N29232 10
D29232 N29232 0 diode
R29233 N29232 N29233 10
D29233 N29233 0 diode
R29234 N29233 N29234 10
D29234 N29234 0 diode
R29235 N29234 N29235 10
D29235 N29235 0 diode
R29236 N29235 N29236 10
D29236 N29236 0 diode
R29237 N29236 N29237 10
D29237 N29237 0 diode
R29238 N29237 N29238 10
D29238 N29238 0 diode
R29239 N29238 N29239 10
D29239 N29239 0 diode
R29240 N29239 N29240 10
D29240 N29240 0 diode
R29241 N29240 N29241 10
D29241 N29241 0 diode
R29242 N29241 N29242 10
D29242 N29242 0 diode
R29243 N29242 N29243 10
D29243 N29243 0 diode
R29244 N29243 N29244 10
D29244 N29244 0 diode
R29245 N29244 N29245 10
D29245 N29245 0 diode
R29246 N29245 N29246 10
D29246 N29246 0 diode
R29247 N29246 N29247 10
D29247 N29247 0 diode
R29248 N29247 N29248 10
D29248 N29248 0 diode
R29249 N29248 N29249 10
D29249 N29249 0 diode
R29250 N29249 N29250 10
D29250 N29250 0 diode
R29251 N29250 N29251 10
D29251 N29251 0 diode
R29252 N29251 N29252 10
D29252 N29252 0 diode
R29253 N29252 N29253 10
D29253 N29253 0 diode
R29254 N29253 N29254 10
D29254 N29254 0 diode
R29255 N29254 N29255 10
D29255 N29255 0 diode
R29256 N29255 N29256 10
D29256 N29256 0 diode
R29257 N29256 N29257 10
D29257 N29257 0 diode
R29258 N29257 N29258 10
D29258 N29258 0 diode
R29259 N29258 N29259 10
D29259 N29259 0 diode
R29260 N29259 N29260 10
D29260 N29260 0 diode
R29261 N29260 N29261 10
D29261 N29261 0 diode
R29262 N29261 N29262 10
D29262 N29262 0 diode
R29263 N29262 N29263 10
D29263 N29263 0 diode
R29264 N29263 N29264 10
D29264 N29264 0 diode
R29265 N29264 N29265 10
D29265 N29265 0 diode
R29266 N29265 N29266 10
D29266 N29266 0 diode
R29267 N29266 N29267 10
D29267 N29267 0 diode
R29268 N29267 N29268 10
D29268 N29268 0 diode
R29269 N29268 N29269 10
D29269 N29269 0 diode
R29270 N29269 N29270 10
D29270 N29270 0 diode
R29271 N29270 N29271 10
D29271 N29271 0 diode
R29272 N29271 N29272 10
D29272 N29272 0 diode
R29273 N29272 N29273 10
D29273 N29273 0 diode
R29274 N29273 N29274 10
D29274 N29274 0 diode
R29275 N29274 N29275 10
D29275 N29275 0 diode
R29276 N29275 N29276 10
D29276 N29276 0 diode
R29277 N29276 N29277 10
D29277 N29277 0 diode
R29278 N29277 N29278 10
D29278 N29278 0 diode
R29279 N29278 N29279 10
D29279 N29279 0 diode
R29280 N29279 N29280 10
D29280 N29280 0 diode
R29281 N29280 N29281 10
D29281 N29281 0 diode
R29282 N29281 N29282 10
D29282 N29282 0 diode
R29283 N29282 N29283 10
D29283 N29283 0 diode
R29284 N29283 N29284 10
D29284 N29284 0 diode
R29285 N29284 N29285 10
D29285 N29285 0 diode
R29286 N29285 N29286 10
D29286 N29286 0 diode
R29287 N29286 N29287 10
D29287 N29287 0 diode
R29288 N29287 N29288 10
D29288 N29288 0 diode
R29289 N29288 N29289 10
D29289 N29289 0 diode
R29290 N29289 N29290 10
D29290 N29290 0 diode
R29291 N29290 N29291 10
D29291 N29291 0 diode
R29292 N29291 N29292 10
D29292 N29292 0 diode
R29293 N29292 N29293 10
D29293 N29293 0 diode
R29294 N29293 N29294 10
D29294 N29294 0 diode
R29295 N29294 N29295 10
D29295 N29295 0 diode
R29296 N29295 N29296 10
D29296 N29296 0 diode
R29297 N29296 N29297 10
D29297 N29297 0 diode
R29298 N29297 N29298 10
D29298 N29298 0 diode
R29299 N29298 N29299 10
D29299 N29299 0 diode
R29300 N29299 N29300 10
D29300 N29300 0 diode
R29301 N29300 N29301 10
D29301 N29301 0 diode
R29302 N29301 N29302 10
D29302 N29302 0 diode
R29303 N29302 N29303 10
D29303 N29303 0 diode
R29304 N29303 N29304 10
D29304 N29304 0 diode
R29305 N29304 N29305 10
D29305 N29305 0 diode
R29306 N29305 N29306 10
D29306 N29306 0 diode
R29307 N29306 N29307 10
D29307 N29307 0 diode
R29308 N29307 N29308 10
D29308 N29308 0 diode
R29309 N29308 N29309 10
D29309 N29309 0 diode
R29310 N29309 N29310 10
D29310 N29310 0 diode
R29311 N29310 N29311 10
D29311 N29311 0 diode
R29312 N29311 N29312 10
D29312 N29312 0 diode
R29313 N29312 N29313 10
D29313 N29313 0 diode
R29314 N29313 N29314 10
D29314 N29314 0 diode
R29315 N29314 N29315 10
D29315 N29315 0 diode
R29316 N29315 N29316 10
D29316 N29316 0 diode
R29317 N29316 N29317 10
D29317 N29317 0 diode
R29318 N29317 N29318 10
D29318 N29318 0 diode
R29319 N29318 N29319 10
D29319 N29319 0 diode
R29320 N29319 N29320 10
D29320 N29320 0 diode
R29321 N29320 N29321 10
D29321 N29321 0 diode
R29322 N29321 N29322 10
D29322 N29322 0 diode
R29323 N29322 N29323 10
D29323 N29323 0 diode
R29324 N29323 N29324 10
D29324 N29324 0 diode
R29325 N29324 N29325 10
D29325 N29325 0 diode
R29326 N29325 N29326 10
D29326 N29326 0 diode
R29327 N29326 N29327 10
D29327 N29327 0 diode
R29328 N29327 N29328 10
D29328 N29328 0 diode
R29329 N29328 N29329 10
D29329 N29329 0 diode
R29330 N29329 N29330 10
D29330 N29330 0 diode
R29331 N29330 N29331 10
D29331 N29331 0 diode
R29332 N29331 N29332 10
D29332 N29332 0 diode
R29333 N29332 N29333 10
D29333 N29333 0 diode
R29334 N29333 N29334 10
D29334 N29334 0 diode
R29335 N29334 N29335 10
D29335 N29335 0 diode
R29336 N29335 N29336 10
D29336 N29336 0 diode
R29337 N29336 N29337 10
D29337 N29337 0 diode
R29338 N29337 N29338 10
D29338 N29338 0 diode
R29339 N29338 N29339 10
D29339 N29339 0 diode
R29340 N29339 N29340 10
D29340 N29340 0 diode
R29341 N29340 N29341 10
D29341 N29341 0 diode
R29342 N29341 N29342 10
D29342 N29342 0 diode
R29343 N29342 N29343 10
D29343 N29343 0 diode
R29344 N29343 N29344 10
D29344 N29344 0 diode
R29345 N29344 N29345 10
D29345 N29345 0 diode
R29346 N29345 N29346 10
D29346 N29346 0 diode
R29347 N29346 N29347 10
D29347 N29347 0 diode
R29348 N29347 N29348 10
D29348 N29348 0 diode
R29349 N29348 N29349 10
D29349 N29349 0 diode
R29350 N29349 N29350 10
D29350 N29350 0 diode
R29351 N29350 N29351 10
D29351 N29351 0 diode
R29352 N29351 N29352 10
D29352 N29352 0 diode
R29353 N29352 N29353 10
D29353 N29353 0 diode
R29354 N29353 N29354 10
D29354 N29354 0 diode
R29355 N29354 N29355 10
D29355 N29355 0 diode
R29356 N29355 N29356 10
D29356 N29356 0 diode
R29357 N29356 N29357 10
D29357 N29357 0 diode
R29358 N29357 N29358 10
D29358 N29358 0 diode
R29359 N29358 N29359 10
D29359 N29359 0 diode
R29360 N29359 N29360 10
D29360 N29360 0 diode
R29361 N29360 N29361 10
D29361 N29361 0 diode
R29362 N29361 N29362 10
D29362 N29362 0 diode
R29363 N29362 N29363 10
D29363 N29363 0 diode
R29364 N29363 N29364 10
D29364 N29364 0 diode
R29365 N29364 N29365 10
D29365 N29365 0 diode
R29366 N29365 N29366 10
D29366 N29366 0 diode
R29367 N29366 N29367 10
D29367 N29367 0 diode
R29368 N29367 N29368 10
D29368 N29368 0 diode
R29369 N29368 N29369 10
D29369 N29369 0 diode
R29370 N29369 N29370 10
D29370 N29370 0 diode
R29371 N29370 N29371 10
D29371 N29371 0 diode
R29372 N29371 N29372 10
D29372 N29372 0 diode
R29373 N29372 N29373 10
D29373 N29373 0 diode
R29374 N29373 N29374 10
D29374 N29374 0 diode
R29375 N29374 N29375 10
D29375 N29375 0 diode
R29376 N29375 N29376 10
D29376 N29376 0 diode
R29377 N29376 N29377 10
D29377 N29377 0 diode
R29378 N29377 N29378 10
D29378 N29378 0 diode
R29379 N29378 N29379 10
D29379 N29379 0 diode
R29380 N29379 N29380 10
D29380 N29380 0 diode
R29381 N29380 N29381 10
D29381 N29381 0 diode
R29382 N29381 N29382 10
D29382 N29382 0 diode
R29383 N29382 N29383 10
D29383 N29383 0 diode
R29384 N29383 N29384 10
D29384 N29384 0 diode
R29385 N29384 N29385 10
D29385 N29385 0 diode
R29386 N29385 N29386 10
D29386 N29386 0 diode
R29387 N29386 N29387 10
D29387 N29387 0 diode
R29388 N29387 N29388 10
D29388 N29388 0 diode
R29389 N29388 N29389 10
D29389 N29389 0 diode
R29390 N29389 N29390 10
D29390 N29390 0 diode
R29391 N29390 N29391 10
D29391 N29391 0 diode
R29392 N29391 N29392 10
D29392 N29392 0 diode
R29393 N29392 N29393 10
D29393 N29393 0 diode
R29394 N29393 N29394 10
D29394 N29394 0 diode
R29395 N29394 N29395 10
D29395 N29395 0 diode
R29396 N29395 N29396 10
D29396 N29396 0 diode
R29397 N29396 N29397 10
D29397 N29397 0 diode
R29398 N29397 N29398 10
D29398 N29398 0 diode
R29399 N29398 N29399 10
D29399 N29399 0 diode
R29400 N29399 N29400 10
D29400 N29400 0 diode
R29401 N29400 N29401 10
D29401 N29401 0 diode
R29402 N29401 N29402 10
D29402 N29402 0 diode
R29403 N29402 N29403 10
D29403 N29403 0 diode
R29404 N29403 N29404 10
D29404 N29404 0 diode
R29405 N29404 N29405 10
D29405 N29405 0 diode
R29406 N29405 N29406 10
D29406 N29406 0 diode
R29407 N29406 N29407 10
D29407 N29407 0 diode
R29408 N29407 N29408 10
D29408 N29408 0 diode
R29409 N29408 N29409 10
D29409 N29409 0 diode
R29410 N29409 N29410 10
D29410 N29410 0 diode
R29411 N29410 N29411 10
D29411 N29411 0 diode
R29412 N29411 N29412 10
D29412 N29412 0 diode
R29413 N29412 N29413 10
D29413 N29413 0 diode
R29414 N29413 N29414 10
D29414 N29414 0 diode
R29415 N29414 N29415 10
D29415 N29415 0 diode
R29416 N29415 N29416 10
D29416 N29416 0 diode
R29417 N29416 N29417 10
D29417 N29417 0 diode
R29418 N29417 N29418 10
D29418 N29418 0 diode
R29419 N29418 N29419 10
D29419 N29419 0 diode
R29420 N29419 N29420 10
D29420 N29420 0 diode
R29421 N29420 N29421 10
D29421 N29421 0 diode
R29422 N29421 N29422 10
D29422 N29422 0 diode
R29423 N29422 N29423 10
D29423 N29423 0 diode
R29424 N29423 N29424 10
D29424 N29424 0 diode
R29425 N29424 N29425 10
D29425 N29425 0 diode
R29426 N29425 N29426 10
D29426 N29426 0 diode
R29427 N29426 N29427 10
D29427 N29427 0 diode
R29428 N29427 N29428 10
D29428 N29428 0 diode
R29429 N29428 N29429 10
D29429 N29429 0 diode
R29430 N29429 N29430 10
D29430 N29430 0 diode
R29431 N29430 N29431 10
D29431 N29431 0 diode
R29432 N29431 N29432 10
D29432 N29432 0 diode
R29433 N29432 N29433 10
D29433 N29433 0 diode
R29434 N29433 N29434 10
D29434 N29434 0 diode
R29435 N29434 N29435 10
D29435 N29435 0 diode
R29436 N29435 N29436 10
D29436 N29436 0 diode
R29437 N29436 N29437 10
D29437 N29437 0 diode
R29438 N29437 N29438 10
D29438 N29438 0 diode
R29439 N29438 N29439 10
D29439 N29439 0 diode
R29440 N29439 N29440 10
D29440 N29440 0 diode
R29441 N29440 N29441 10
D29441 N29441 0 diode
R29442 N29441 N29442 10
D29442 N29442 0 diode
R29443 N29442 N29443 10
D29443 N29443 0 diode
R29444 N29443 N29444 10
D29444 N29444 0 diode
R29445 N29444 N29445 10
D29445 N29445 0 diode
R29446 N29445 N29446 10
D29446 N29446 0 diode
R29447 N29446 N29447 10
D29447 N29447 0 diode
R29448 N29447 N29448 10
D29448 N29448 0 diode
R29449 N29448 N29449 10
D29449 N29449 0 diode
R29450 N29449 N29450 10
D29450 N29450 0 diode
R29451 N29450 N29451 10
D29451 N29451 0 diode
R29452 N29451 N29452 10
D29452 N29452 0 diode
R29453 N29452 N29453 10
D29453 N29453 0 diode
R29454 N29453 N29454 10
D29454 N29454 0 diode
R29455 N29454 N29455 10
D29455 N29455 0 diode
R29456 N29455 N29456 10
D29456 N29456 0 diode
R29457 N29456 N29457 10
D29457 N29457 0 diode
R29458 N29457 N29458 10
D29458 N29458 0 diode
R29459 N29458 N29459 10
D29459 N29459 0 diode
R29460 N29459 N29460 10
D29460 N29460 0 diode
R29461 N29460 N29461 10
D29461 N29461 0 diode
R29462 N29461 N29462 10
D29462 N29462 0 diode
R29463 N29462 N29463 10
D29463 N29463 0 diode
R29464 N29463 N29464 10
D29464 N29464 0 diode
R29465 N29464 N29465 10
D29465 N29465 0 diode
R29466 N29465 N29466 10
D29466 N29466 0 diode
R29467 N29466 N29467 10
D29467 N29467 0 diode
R29468 N29467 N29468 10
D29468 N29468 0 diode
R29469 N29468 N29469 10
D29469 N29469 0 diode
R29470 N29469 N29470 10
D29470 N29470 0 diode
R29471 N29470 N29471 10
D29471 N29471 0 diode
R29472 N29471 N29472 10
D29472 N29472 0 diode
R29473 N29472 N29473 10
D29473 N29473 0 diode
R29474 N29473 N29474 10
D29474 N29474 0 diode
R29475 N29474 N29475 10
D29475 N29475 0 diode
R29476 N29475 N29476 10
D29476 N29476 0 diode
R29477 N29476 N29477 10
D29477 N29477 0 diode
R29478 N29477 N29478 10
D29478 N29478 0 diode
R29479 N29478 N29479 10
D29479 N29479 0 diode
R29480 N29479 N29480 10
D29480 N29480 0 diode
R29481 N29480 N29481 10
D29481 N29481 0 diode
R29482 N29481 N29482 10
D29482 N29482 0 diode
R29483 N29482 N29483 10
D29483 N29483 0 diode
R29484 N29483 N29484 10
D29484 N29484 0 diode
R29485 N29484 N29485 10
D29485 N29485 0 diode
R29486 N29485 N29486 10
D29486 N29486 0 diode
R29487 N29486 N29487 10
D29487 N29487 0 diode
R29488 N29487 N29488 10
D29488 N29488 0 diode
R29489 N29488 N29489 10
D29489 N29489 0 diode
R29490 N29489 N29490 10
D29490 N29490 0 diode
R29491 N29490 N29491 10
D29491 N29491 0 diode
R29492 N29491 N29492 10
D29492 N29492 0 diode
R29493 N29492 N29493 10
D29493 N29493 0 diode
R29494 N29493 N29494 10
D29494 N29494 0 diode
R29495 N29494 N29495 10
D29495 N29495 0 diode
R29496 N29495 N29496 10
D29496 N29496 0 diode
R29497 N29496 N29497 10
D29497 N29497 0 diode
R29498 N29497 N29498 10
D29498 N29498 0 diode
R29499 N29498 N29499 10
D29499 N29499 0 diode
R29500 N29499 N29500 10
D29500 N29500 0 diode
R29501 N29500 N29501 10
D29501 N29501 0 diode
R29502 N29501 N29502 10
D29502 N29502 0 diode
R29503 N29502 N29503 10
D29503 N29503 0 diode
R29504 N29503 N29504 10
D29504 N29504 0 diode
R29505 N29504 N29505 10
D29505 N29505 0 diode
R29506 N29505 N29506 10
D29506 N29506 0 diode
R29507 N29506 N29507 10
D29507 N29507 0 diode
R29508 N29507 N29508 10
D29508 N29508 0 diode
R29509 N29508 N29509 10
D29509 N29509 0 diode
R29510 N29509 N29510 10
D29510 N29510 0 diode
R29511 N29510 N29511 10
D29511 N29511 0 diode
R29512 N29511 N29512 10
D29512 N29512 0 diode
R29513 N29512 N29513 10
D29513 N29513 0 diode
R29514 N29513 N29514 10
D29514 N29514 0 diode
R29515 N29514 N29515 10
D29515 N29515 0 diode
R29516 N29515 N29516 10
D29516 N29516 0 diode
R29517 N29516 N29517 10
D29517 N29517 0 diode
R29518 N29517 N29518 10
D29518 N29518 0 diode
R29519 N29518 N29519 10
D29519 N29519 0 diode
R29520 N29519 N29520 10
D29520 N29520 0 diode
R29521 N29520 N29521 10
D29521 N29521 0 diode
R29522 N29521 N29522 10
D29522 N29522 0 diode
R29523 N29522 N29523 10
D29523 N29523 0 diode
R29524 N29523 N29524 10
D29524 N29524 0 diode
R29525 N29524 N29525 10
D29525 N29525 0 diode
R29526 N29525 N29526 10
D29526 N29526 0 diode
R29527 N29526 N29527 10
D29527 N29527 0 diode
R29528 N29527 N29528 10
D29528 N29528 0 diode
R29529 N29528 N29529 10
D29529 N29529 0 diode
R29530 N29529 N29530 10
D29530 N29530 0 diode
R29531 N29530 N29531 10
D29531 N29531 0 diode
R29532 N29531 N29532 10
D29532 N29532 0 diode
R29533 N29532 N29533 10
D29533 N29533 0 diode
R29534 N29533 N29534 10
D29534 N29534 0 diode
R29535 N29534 N29535 10
D29535 N29535 0 diode
R29536 N29535 N29536 10
D29536 N29536 0 diode
R29537 N29536 N29537 10
D29537 N29537 0 diode
R29538 N29537 N29538 10
D29538 N29538 0 diode
R29539 N29538 N29539 10
D29539 N29539 0 diode
R29540 N29539 N29540 10
D29540 N29540 0 diode
R29541 N29540 N29541 10
D29541 N29541 0 diode
R29542 N29541 N29542 10
D29542 N29542 0 diode
R29543 N29542 N29543 10
D29543 N29543 0 diode
R29544 N29543 N29544 10
D29544 N29544 0 diode
R29545 N29544 N29545 10
D29545 N29545 0 diode
R29546 N29545 N29546 10
D29546 N29546 0 diode
R29547 N29546 N29547 10
D29547 N29547 0 diode
R29548 N29547 N29548 10
D29548 N29548 0 diode
R29549 N29548 N29549 10
D29549 N29549 0 diode
R29550 N29549 N29550 10
D29550 N29550 0 diode
R29551 N29550 N29551 10
D29551 N29551 0 diode
R29552 N29551 N29552 10
D29552 N29552 0 diode
R29553 N29552 N29553 10
D29553 N29553 0 diode
R29554 N29553 N29554 10
D29554 N29554 0 diode
R29555 N29554 N29555 10
D29555 N29555 0 diode
R29556 N29555 N29556 10
D29556 N29556 0 diode
R29557 N29556 N29557 10
D29557 N29557 0 diode
R29558 N29557 N29558 10
D29558 N29558 0 diode
R29559 N29558 N29559 10
D29559 N29559 0 diode
R29560 N29559 N29560 10
D29560 N29560 0 diode
R29561 N29560 N29561 10
D29561 N29561 0 diode
R29562 N29561 N29562 10
D29562 N29562 0 diode
R29563 N29562 N29563 10
D29563 N29563 0 diode
R29564 N29563 N29564 10
D29564 N29564 0 diode
R29565 N29564 N29565 10
D29565 N29565 0 diode
R29566 N29565 N29566 10
D29566 N29566 0 diode
R29567 N29566 N29567 10
D29567 N29567 0 diode
R29568 N29567 N29568 10
D29568 N29568 0 diode
R29569 N29568 N29569 10
D29569 N29569 0 diode
R29570 N29569 N29570 10
D29570 N29570 0 diode
R29571 N29570 N29571 10
D29571 N29571 0 diode
R29572 N29571 N29572 10
D29572 N29572 0 diode
R29573 N29572 N29573 10
D29573 N29573 0 diode
R29574 N29573 N29574 10
D29574 N29574 0 diode
R29575 N29574 N29575 10
D29575 N29575 0 diode
R29576 N29575 N29576 10
D29576 N29576 0 diode
R29577 N29576 N29577 10
D29577 N29577 0 diode
R29578 N29577 N29578 10
D29578 N29578 0 diode
R29579 N29578 N29579 10
D29579 N29579 0 diode
R29580 N29579 N29580 10
D29580 N29580 0 diode
R29581 N29580 N29581 10
D29581 N29581 0 diode
R29582 N29581 N29582 10
D29582 N29582 0 diode
R29583 N29582 N29583 10
D29583 N29583 0 diode
R29584 N29583 N29584 10
D29584 N29584 0 diode
R29585 N29584 N29585 10
D29585 N29585 0 diode
R29586 N29585 N29586 10
D29586 N29586 0 diode
R29587 N29586 N29587 10
D29587 N29587 0 diode
R29588 N29587 N29588 10
D29588 N29588 0 diode
R29589 N29588 N29589 10
D29589 N29589 0 diode
R29590 N29589 N29590 10
D29590 N29590 0 diode
R29591 N29590 N29591 10
D29591 N29591 0 diode
R29592 N29591 N29592 10
D29592 N29592 0 diode
R29593 N29592 N29593 10
D29593 N29593 0 diode
R29594 N29593 N29594 10
D29594 N29594 0 diode
R29595 N29594 N29595 10
D29595 N29595 0 diode
R29596 N29595 N29596 10
D29596 N29596 0 diode
R29597 N29596 N29597 10
D29597 N29597 0 diode
R29598 N29597 N29598 10
D29598 N29598 0 diode
R29599 N29598 N29599 10
D29599 N29599 0 diode
R29600 N29599 N29600 10
D29600 N29600 0 diode
R29601 N29600 N29601 10
D29601 N29601 0 diode
R29602 N29601 N29602 10
D29602 N29602 0 diode
R29603 N29602 N29603 10
D29603 N29603 0 diode
R29604 N29603 N29604 10
D29604 N29604 0 diode
R29605 N29604 N29605 10
D29605 N29605 0 diode
R29606 N29605 N29606 10
D29606 N29606 0 diode
R29607 N29606 N29607 10
D29607 N29607 0 diode
R29608 N29607 N29608 10
D29608 N29608 0 diode
R29609 N29608 N29609 10
D29609 N29609 0 diode
R29610 N29609 N29610 10
D29610 N29610 0 diode
R29611 N29610 N29611 10
D29611 N29611 0 diode
R29612 N29611 N29612 10
D29612 N29612 0 diode
R29613 N29612 N29613 10
D29613 N29613 0 diode
R29614 N29613 N29614 10
D29614 N29614 0 diode
R29615 N29614 N29615 10
D29615 N29615 0 diode
R29616 N29615 N29616 10
D29616 N29616 0 diode
R29617 N29616 N29617 10
D29617 N29617 0 diode
R29618 N29617 N29618 10
D29618 N29618 0 diode
R29619 N29618 N29619 10
D29619 N29619 0 diode
R29620 N29619 N29620 10
D29620 N29620 0 diode
R29621 N29620 N29621 10
D29621 N29621 0 diode
R29622 N29621 N29622 10
D29622 N29622 0 diode
R29623 N29622 N29623 10
D29623 N29623 0 diode
R29624 N29623 N29624 10
D29624 N29624 0 diode
R29625 N29624 N29625 10
D29625 N29625 0 diode
R29626 N29625 N29626 10
D29626 N29626 0 diode
R29627 N29626 N29627 10
D29627 N29627 0 diode
R29628 N29627 N29628 10
D29628 N29628 0 diode
R29629 N29628 N29629 10
D29629 N29629 0 diode
R29630 N29629 N29630 10
D29630 N29630 0 diode
R29631 N29630 N29631 10
D29631 N29631 0 diode
R29632 N29631 N29632 10
D29632 N29632 0 diode
R29633 N29632 N29633 10
D29633 N29633 0 diode
R29634 N29633 N29634 10
D29634 N29634 0 diode
R29635 N29634 N29635 10
D29635 N29635 0 diode
R29636 N29635 N29636 10
D29636 N29636 0 diode
R29637 N29636 N29637 10
D29637 N29637 0 diode
R29638 N29637 N29638 10
D29638 N29638 0 diode
R29639 N29638 N29639 10
D29639 N29639 0 diode
R29640 N29639 N29640 10
D29640 N29640 0 diode
R29641 N29640 N29641 10
D29641 N29641 0 diode
R29642 N29641 N29642 10
D29642 N29642 0 diode
R29643 N29642 N29643 10
D29643 N29643 0 diode
R29644 N29643 N29644 10
D29644 N29644 0 diode
R29645 N29644 N29645 10
D29645 N29645 0 diode
R29646 N29645 N29646 10
D29646 N29646 0 diode
R29647 N29646 N29647 10
D29647 N29647 0 diode
R29648 N29647 N29648 10
D29648 N29648 0 diode
R29649 N29648 N29649 10
D29649 N29649 0 diode
R29650 N29649 N29650 10
D29650 N29650 0 diode
R29651 N29650 N29651 10
D29651 N29651 0 diode
R29652 N29651 N29652 10
D29652 N29652 0 diode
R29653 N29652 N29653 10
D29653 N29653 0 diode
R29654 N29653 N29654 10
D29654 N29654 0 diode
R29655 N29654 N29655 10
D29655 N29655 0 diode
R29656 N29655 N29656 10
D29656 N29656 0 diode
R29657 N29656 N29657 10
D29657 N29657 0 diode
R29658 N29657 N29658 10
D29658 N29658 0 diode
R29659 N29658 N29659 10
D29659 N29659 0 diode
R29660 N29659 N29660 10
D29660 N29660 0 diode
R29661 N29660 N29661 10
D29661 N29661 0 diode
R29662 N29661 N29662 10
D29662 N29662 0 diode
R29663 N29662 N29663 10
D29663 N29663 0 diode
R29664 N29663 N29664 10
D29664 N29664 0 diode
R29665 N29664 N29665 10
D29665 N29665 0 diode
R29666 N29665 N29666 10
D29666 N29666 0 diode
R29667 N29666 N29667 10
D29667 N29667 0 diode
R29668 N29667 N29668 10
D29668 N29668 0 diode
R29669 N29668 N29669 10
D29669 N29669 0 diode
R29670 N29669 N29670 10
D29670 N29670 0 diode
R29671 N29670 N29671 10
D29671 N29671 0 diode
R29672 N29671 N29672 10
D29672 N29672 0 diode
R29673 N29672 N29673 10
D29673 N29673 0 diode
R29674 N29673 N29674 10
D29674 N29674 0 diode
R29675 N29674 N29675 10
D29675 N29675 0 diode
R29676 N29675 N29676 10
D29676 N29676 0 diode
R29677 N29676 N29677 10
D29677 N29677 0 diode
R29678 N29677 N29678 10
D29678 N29678 0 diode
R29679 N29678 N29679 10
D29679 N29679 0 diode
R29680 N29679 N29680 10
D29680 N29680 0 diode
R29681 N29680 N29681 10
D29681 N29681 0 diode
R29682 N29681 N29682 10
D29682 N29682 0 diode
R29683 N29682 N29683 10
D29683 N29683 0 diode
R29684 N29683 N29684 10
D29684 N29684 0 diode
R29685 N29684 N29685 10
D29685 N29685 0 diode
R29686 N29685 N29686 10
D29686 N29686 0 diode
R29687 N29686 N29687 10
D29687 N29687 0 diode
R29688 N29687 N29688 10
D29688 N29688 0 diode
R29689 N29688 N29689 10
D29689 N29689 0 diode
R29690 N29689 N29690 10
D29690 N29690 0 diode
R29691 N29690 N29691 10
D29691 N29691 0 diode
R29692 N29691 N29692 10
D29692 N29692 0 diode
R29693 N29692 N29693 10
D29693 N29693 0 diode
R29694 N29693 N29694 10
D29694 N29694 0 diode
R29695 N29694 N29695 10
D29695 N29695 0 diode
R29696 N29695 N29696 10
D29696 N29696 0 diode
R29697 N29696 N29697 10
D29697 N29697 0 diode
R29698 N29697 N29698 10
D29698 N29698 0 diode
R29699 N29698 N29699 10
D29699 N29699 0 diode
R29700 N29699 N29700 10
D29700 N29700 0 diode
R29701 N29700 N29701 10
D29701 N29701 0 diode
R29702 N29701 N29702 10
D29702 N29702 0 diode
R29703 N29702 N29703 10
D29703 N29703 0 diode
R29704 N29703 N29704 10
D29704 N29704 0 diode
R29705 N29704 N29705 10
D29705 N29705 0 diode
R29706 N29705 N29706 10
D29706 N29706 0 diode
R29707 N29706 N29707 10
D29707 N29707 0 diode
R29708 N29707 N29708 10
D29708 N29708 0 diode
R29709 N29708 N29709 10
D29709 N29709 0 diode
R29710 N29709 N29710 10
D29710 N29710 0 diode
R29711 N29710 N29711 10
D29711 N29711 0 diode
R29712 N29711 N29712 10
D29712 N29712 0 diode
R29713 N29712 N29713 10
D29713 N29713 0 diode
R29714 N29713 N29714 10
D29714 N29714 0 diode
R29715 N29714 N29715 10
D29715 N29715 0 diode
R29716 N29715 N29716 10
D29716 N29716 0 diode
R29717 N29716 N29717 10
D29717 N29717 0 diode
R29718 N29717 N29718 10
D29718 N29718 0 diode
R29719 N29718 N29719 10
D29719 N29719 0 diode
R29720 N29719 N29720 10
D29720 N29720 0 diode
R29721 N29720 N29721 10
D29721 N29721 0 diode
R29722 N29721 N29722 10
D29722 N29722 0 diode
R29723 N29722 N29723 10
D29723 N29723 0 diode
R29724 N29723 N29724 10
D29724 N29724 0 diode
R29725 N29724 N29725 10
D29725 N29725 0 diode
R29726 N29725 N29726 10
D29726 N29726 0 diode
R29727 N29726 N29727 10
D29727 N29727 0 diode
R29728 N29727 N29728 10
D29728 N29728 0 diode
R29729 N29728 N29729 10
D29729 N29729 0 diode
R29730 N29729 N29730 10
D29730 N29730 0 diode
R29731 N29730 N29731 10
D29731 N29731 0 diode
R29732 N29731 N29732 10
D29732 N29732 0 diode
R29733 N29732 N29733 10
D29733 N29733 0 diode
R29734 N29733 N29734 10
D29734 N29734 0 diode
R29735 N29734 N29735 10
D29735 N29735 0 diode
R29736 N29735 N29736 10
D29736 N29736 0 diode
R29737 N29736 N29737 10
D29737 N29737 0 diode
R29738 N29737 N29738 10
D29738 N29738 0 diode
R29739 N29738 N29739 10
D29739 N29739 0 diode
R29740 N29739 N29740 10
D29740 N29740 0 diode
R29741 N29740 N29741 10
D29741 N29741 0 diode
R29742 N29741 N29742 10
D29742 N29742 0 diode
R29743 N29742 N29743 10
D29743 N29743 0 diode
R29744 N29743 N29744 10
D29744 N29744 0 diode
R29745 N29744 N29745 10
D29745 N29745 0 diode
R29746 N29745 N29746 10
D29746 N29746 0 diode
R29747 N29746 N29747 10
D29747 N29747 0 diode
R29748 N29747 N29748 10
D29748 N29748 0 diode
R29749 N29748 N29749 10
D29749 N29749 0 diode
R29750 N29749 N29750 10
D29750 N29750 0 diode
R29751 N29750 N29751 10
D29751 N29751 0 diode
R29752 N29751 N29752 10
D29752 N29752 0 diode
R29753 N29752 N29753 10
D29753 N29753 0 diode
R29754 N29753 N29754 10
D29754 N29754 0 diode
R29755 N29754 N29755 10
D29755 N29755 0 diode
R29756 N29755 N29756 10
D29756 N29756 0 diode
R29757 N29756 N29757 10
D29757 N29757 0 diode
R29758 N29757 N29758 10
D29758 N29758 0 diode
R29759 N29758 N29759 10
D29759 N29759 0 diode
R29760 N29759 N29760 10
D29760 N29760 0 diode
R29761 N29760 N29761 10
D29761 N29761 0 diode
R29762 N29761 N29762 10
D29762 N29762 0 diode
R29763 N29762 N29763 10
D29763 N29763 0 diode
R29764 N29763 N29764 10
D29764 N29764 0 diode
R29765 N29764 N29765 10
D29765 N29765 0 diode
R29766 N29765 N29766 10
D29766 N29766 0 diode
R29767 N29766 N29767 10
D29767 N29767 0 diode
R29768 N29767 N29768 10
D29768 N29768 0 diode
R29769 N29768 N29769 10
D29769 N29769 0 diode
R29770 N29769 N29770 10
D29770 N29770 0 diode
R29771 N29770 N29771 10
D29771 N29771 0 diode
R29772 N29771 N29772 10
D29772 N29772 0 diode
R29773 N29772 N29773 10
D29773 N29773 0 diode
R29774 N29773 N29774 10
D29774 N29774 0 diode
R29775 N29774 N29775 10
D29775 N29775 0 diode
R29776 N29775 N29776 10
D29776 N29776 0 diode
R29777 N29776 N29777 10
D29777 N29777 0 diode
R29778 N29777 N29778 10
D29778 N29778 0 diode
R29779 N29778 N29779 10
D29779 N29779 0 diode
R29780 N29779 N29780 10
D29780 N29780 0 diode
R29781 N29780 N29781 10
D29781 N29781 0 diode
R29782 N29781 N29782 10
D29782 N29782 0 diode
R29783 N29782 N29783 10
D29783 N29783 0 diode
R29784 N29783 N29784 10
D29784 N29784 0 diode
R29785 N29784 N29785 10
D29785 N29785 0 diode
R29786 N29785 N29786 10
D29786 N29786 0 diode
R29787 N29786 N29787 10
D29787 N29787 0 diode
R29788 N29787 N29788 10
D29788 N29788 0 diode
R29789 N29788 N29789 10
D29789 N29789 0 diode
R29790 N29789 N29790 10
D29790 N29790 0 diode
R29791 N29790 N29791 10
D29791 N29791 0 diode
R29792 N29791 N29792 10
D29792 N29792 0 diode
R29793 N29792 N29793 10
D29793 N29793 0 diode
R29794 N29793 N29794 10
D29794 N29794 0 diode
R29795 N29794 N29795 10
D29795 N29795 0 diode
R29796 N29795 N29796 10
D29796 N29796 0 diode
R29797 N29796 N29797 10
D29797 N29797 0 diode
R29798 N29797 N29798 10
D29798 N29798 0 diode
R29799 N29798 N29799 10
D29799 N29799 0 diode
R29800 N29799 N29800 10
D29800 N29800 0 diode
R29801 N29800 N29801 10
D29801 N29801 0 diode
R29802 N29801 N29802 10
D29802 N29802 0 diode
R29803 N29802 N29803 10
D29803 N29803 0 diode
R29804 N29803 N29804 10
D29804 N29804 0 diode
R29805 N29804 N29805 10
D29805 N29805 0 diode
R29806 N29805 N29806 10
D29806 N29806 0 diode
R29807 N29806 N29807 10
D29807 N29807 0 diode
R29808 N29807 N29808 10
D29808 N29808 0 diode
R29809 N29808 N29809 10
D29809 N29809 0 diode
R29810 N29809 N29810 10
D29810 N29810 0 diode
R29811 N29810 N29811 10
D29811 N29811 0 diode
R29812 N29811 N29812 10
D29812 N29812 0 diode
R29813 N29812 N29813 10
D29813 N29813 0 diode
R29814 N29813 N29814 10
D29814 N29814 0 diode
R29815 N29814 N29815 10
D29815 N29815 0 diode
R29816 N29815 N29816 10
D29816 N29816 0 diode
R29817 N29816 N29817 10
D29817 N29817 0 diode
R29818 N29817 N29818 10
D29818 N29818 0 diode
R29819 N29818 N29819 10
D29819 N29819 0 diode
R29820 N29819 N29820 10
D29820 N29820 0 diode
R29821 N29820 N29821 10
D29821 N29821 0 diode
R29822 N29821 N29822 10
D29822 N29822 0 diode
R29823 N29822 N29823 10
D29823 N29823 0 diode
R29824 N29823 N29824 10
D29824 N29824 0 diode
R29825 N29824 N29825 10
D29825 N29825 0 diode
R29826 N29825 N29826 10
D29826 N29826 0 diode
R29827 N29826 N29827 10
D29827 N29827 0 diode
R29828 N29827 N29828 10
D29828 N29828 0 diode
R29829 N29828 N29829 10
D29829 N29829 0 diode
R29830 N29829 N29830 10
D29830 N29830 0 diode
R29831 N29830 N29831 10
D29831 N29831 0 diode
R29832 N29831 N29832 10
D29832 N29832 0 diode
R29833 N29832 N29833 10
D29833 N29833 0 diode
R29834 N29833 N29834 10
D29834 N29834 0 diode
R29835 N29834 N29835 10
D29835 N29835 0 diode
R29836 N29835 N29836 10
D29836 N29836 0 diode
R29837 N29836 N29837 10
D29837 N29837 0 diode
R29838 N29837 N29838 10
D29838 N29838 0 diode
R29839 N29838 N29839 10
D29839 N29839 0 diode
R29840 N29839 N29840 10
D29840 N29840 0 diode
R29841 N29840 N29841 10
D29841 N29841 0 diode
R29842 N29841 N29842 10
D29842 N29842 0 diode
R29843 N29842 N29843 10
D29843 N29843 0 diode
R29844 N29843 N29844 10
D29844 N29844 0 diode
R29845 N29844 N29845 10
D29845 N29845 0 diode
R29846 N29845 N29846 10
D29846 N29846 0 diode
R29847 N29846 N29847 10
D29847 N29847 0 diode
R29848 N29847 N29848 10
D29848 N29848 0 diode
R29849 N29848 N29849 10
D29849 N29849 0 diode
R29850 N29849 N29850 10
D29850 N29850 0 diode
R29851 N29850 N29851 10
D29851 N29851 0 diode
R29852 N29851 N29852 10
D29852 N29852 0 diode
R29853 N29852 N29853 10
D29853 N29853 0 diode
R29854 N29853 N29854 10
D29854 N29854 0 diode
R29855 N29854 N29855 10
D29855 N29855 0 diode
R29856 N29855 N29856 10
D29856 N29856 0 diode
R29857 N29856 N29857 10
D29857 N29857 0 diode
R29858 N29857 N29858 10
D29858 N29858 0 diode
R29859 N29858 N29859 10
D29859 N29859 0 diode
R29860 N29859 N29860 10
D29860 N29860 0 diode
R29861 N29860 N29861 10
D29861 N29861 0 diode
R29862 N29861 N29862 10
D29862 N29862 0 diode
R29863 N29862 N29863 10
D29863 N29863 0 diode
R29864 N29863 N29864 10
D29864 N29864 0 diode
R29865 N29864 N29865 10
D29865 N29865 0 diode
R29866 N29865 N29866 10
D29866 N29866 0 diode
R29867 N29866 N29867 10
D29867 N29867 0 diode
R29868 N29867 N29868 10
D29868 N29868 0 diode
R29869 N29868 N29869 10
D29869 N29869 0 diode
R29870 N29869 N29870 10
D29870 N29870 0 diode
R29871 N29870 N29871 10
D29871 N29871 0 diode
R29872 N29871 N29872 10
D29872 N29872 0 diode
R29873 N29872 N29873 10
D29873 N29873 0 diode
R29874 N29873 N29874 10
D29874 N29874 0 diode
R29875 N29874 N29875 10
D29875 N29875 0 diode
R29876 N29875 N29876 10
D29876 N29876 0 diode
R29877 N29876 N29877 10
D29877 N29877 0 diode
R29878 N29877 N29878 10
D29878 N29878 0 diode
R29879 N29878 N29879 10
D29879 N29879 0 diode
R29880 N29879 N29880 10
D29880 N29880 0 diode
R29881 N29880 N29881 10
D29881 N29881 0 diode
R29882 N29881 N29882 10
D29882 N29882 0 diode
R29883 N29882 N29883 10
D29883 N29883 0 diode
R29884 N29883 N29884 10
D29884 N29884 0 diode
R29885 N29884 N29885 10
D29885 N29885 0 diode
R29886 N29885 N29886 10
D29886 N29886 0 diode
R29887 N29886 N29887 10
D29887 N29887 0 diode
R29888 N29887 N29888 10
D29888 N29888 0 diode
R29889 N29888 N29889 10
D29889 N29889 0 diode
R29890 N29889 N29890 10
D29890 N29890 0 diode
R29891 N29890 N29891 10
D29891 N29891 0 diode
R29892 N29891 N29892 10
D29892 N29892 0 diode
R29893 N29892 N29893 10
D29893 N29893 0 diode
R29894 N29893 N29894 10
D29894 N29894 0 diode
R29895 N29894 N29895 10
D29895 N29895 0 diode
R29896 N29895 N29896 10
D29896 N29896 0 diode
R29897 N29896 N29897 10
D29897 N29897 0 diode
R29898 N29897 N29898 10
D29898 N29898 0 diode
R29899 N29898 N29899 10
D29899 N29899 0 diode
R29900 N29899 N29900 10
D29900 N29900 0 diode
R29901 N29900 N29901 10
D29901 N29901 0 diode
R29902 N29901 N29902 10
D29902 N29902 0 diode
R29903 N29902 N29903 10
D29903 N29903 0 diode
R29904 N29903 N29904 10
D29904 N29904 0 diode
R29905 N29904 N29905 10
D29905 N29905 0 diode
R29906 N29905 N29906 10
D29906 N29906 0 diode
R29907 N29906 N29907 10
D29907 N29907 0 diode
R29908 N29907 N29908 10
D29908 N29908 0 diode
R29909 N29908 N29909 10
D29909 N29909 0 diode
R29910 N29909 N29910 10
D29910 N29910 0 diode
R29911 N29910 N29911 10
D29911 N29911 0 diode
R29912 N29911 N29912 10
D29912 N29912 0 diode
R29913 N29912 N29913 10
D29913 N29913 0 diode
R29914 N29913 N29914 10
D29914 N29914 0 diode
R29915 N29914 N29915 10
D29915 N29915 0 diode
R29916 N29915 N29916 10
D29916 N29916 0 diode
R29917 N29916 N29917 10
D29917 N29917 0 diode
R29918 N29917 N29918 10
D29918 N29918 0 diode
R29919 N29918 N29919 10
D29919 N29919 0 diode
R29920 N29919 N29920 10
D29920 N29920 0 diode
R29921 N29920 N29921 10
D29921 N29921 0 diode
R29922 N29921 N29922 10
D29922 N29922 0 diode
R29923 N29922 N29923 10
D29923 N29923 0 diode
R29924 N29923 N29924 10
D29924 N29924 0 diode
R29925 N29924 N29925 10
D29925 N29925 0 diode
R29926 N29925 N29926 10
D29926 N29926 0 diode
R29927 N29926 N29927 10
D29927 N29927 0 diode
R29928 N29927 N29928 10
D29928 N29928 0 diode
R29929 N29928 N29929 10
D29929 N29929 0 diode
R29930 N29929 N29930 10
D29930 N29930 0 diode
R29931 N29930 N29931 10
D29931 N29931 0 diode
R29932 N29931 N29932 10
D29932 N29932 0 diode
R29933 N29932 N29933 10
D29933 N29933 0 diode
R29934 N29933 N29934 10
D29934 N29934 0 diode
R29935 N29934 N29935 10
D29935 N29935 0 diode
R29936 N29935 N29936 10
D29936 N29936 0 diode
R29937 N29936 N29937 10
D29937 N29937 0 diode
R29938 N29937 N29938 10
D29938 N29938 0 diode
R29939 N29938 N29939 10
D29939 N29939 0 diode
R29940 N29939 N29940 10
D29940 N29940 0 diode
R29941 N29940 N29941 10
D29941 N29941 0 diode
R29942 N29941 N29942 10
D29942 N29942 0 diode
R29943 N29942 N29943 10
D29943 N29943 0 diode
R29944 N29943 N29944 10
D29944 N29944 0 diode
R29945 N29944 N29945 10
D29945 N29945 0 diode
R29946 N29945 N29946 10
D29946 N29946 0 diode
R29947 N29946 N29947 10
D29947 N29947 0 diode
R29948 N29947 N29948 10
D29948 N29948 0 diode
R29949 N29948 N29949 10
D29949 N29949 0 diode
R29950 N29949 N29950 10
D29950 N29950 0 diode
R29951 N29950 N29951 10
D29951 N29951 0 diode
R29952 N29951 N29952 10
D29952 N29952 0 diode
R29953 N29952 N29953 10
D29953 N29953 0 diode
R29954 N29953 N29954 10
D29954 N29954 0 diode
R29955 N29954 N29955 10
D29955 N29955 0 diode
R29956 N29955 N29956 10
D29956 N29956 0 diode
R29957 N29956 N29957 10
D29957 N29957 0 diode
R29958 N29957 N29958 10
D29958 N29958 0 diode
R29959 N29958 N29959 10
D29959 N29959 0 diode
R29960 N29959 N29960 10
D29960 N29960 0 diode
R29961 N29960 N29961 10
D29961 N29961 0 diode
R29962 N29961 N29962 10
D29962 N29962 0 diode
R29963 N29962 N29963 10
D29963 N29963 0 diode
R29964 N29963 N29964 10
D29964 N29964 0 diode
R29965 N29964 N29965 10
D29965 N29965 0 diode
R29966 N29965 N29966 10
D29966 N29966 0 diode
R29967 N29966 N29967 10
D29967 N29967 0 diode
R29968 N29967 N29968 10
D29968 N29968 0 diode
R29969 N29968 N29969 10
D29969 N29969 0 diode
R29970 N29969 N29970 10
D29970 N29970 0 diode
R29971 N29970 N29971 10
D29971 N29971 0 diode
R29972 N29971 N29972 10
D29972 N29972 0 diode
R29973 N29972 N29973 10
D29973 N29973 0 diode
R29974 N29973 N29974 10
D29974 N29974 0 diode
R29975 N29974 N29975 10
D29975 N29975 0 diode
R29976 N29975 N29976 10
D29976 N29976 0 diode
R29977 N29976 N29977 10
D29977 N29977 0 diode
R29978 N29977 N29978 10
D29978 N29978 0 diode
R29979 N29978 N29979 10
D29979 N29979 0 diode
R29980 N29979 N29980 10
D29980 N29980 0 diode
R29981 N29980 N29981 10
D29981 N29981 0 diode
R29982 N29981 N29982 10
D29982 N29982 0 diode
R29983 N29982 N29983 10
D29983 N29983 0 diode
R29984 N29983 N29984 10
D29984 N29984 0 diode
R29985 N29984 N29985 10
D29985 N29985 0 diode
R29986 N29985 N29986 10
D29986 N29986 0 diode
R29987 N29986 N29987 10
D29987 N29987 0 diode
R29988 N29987 N29988 10
D29988 N29988 0 diode
R29989 N29988 N29989 10
D29989 N29989 0 diode
R29990 N29989 N29990 10
D29990 N29990 0 diode
R29991 N29990 N29991 10
D29991 N29991 0 diode
R29992 N29991 N29992 10
D29992 N29992 0 diode
R29993 N29992 N29993 10
D29993 N29993 0 diode
R29994 N29993 N29994 10
D29994 N29994 0 diode
R29995 N29994 N29995 10
D29995 N29995 0 diode
R29996 N29995 N29996 10
D29996 N29996 0 diode
R29997 N29996 N29997 10
D29997 N29997 0 diode
R29998 N29997 N29998 10
D29998 N29998 0 diode
R29999 N29998 N29999 10
D29999 N29999 0 diode
R30000 N29999 N30000 10
D30000 N30000 0 diode
R30001 N30000 N30001 10
D30001 N30001 0 diode
R30002 N30001 N30002 10
D30002 N30002 0 diode
R30003 N30002 N30003 10
D30003 N30003 0 diode
R30004 N30003 N30004 10
D30004 N30004 0 diode
R30005 N30004 N30005 10
D30005 N30005 0 diode
R30006 N30005 N30006 10
D30006 N30006 0 diode
R30007 N30006 N30007 10
D30007 N30007 0 diode
R30008 N30007 N30008 10
D30008 N30008 0 diode
R30009 N30008 N30009 10
D30009 N30009 0 diode
R30010 N30009 N30010 10
D30010 N30010 0 diode
R30011 N30010 N30011 10
D30011 N30011 0 diode
R30012 N30011 N30012 10
D30012 N30012 0 diode
R30013 N30012 N30013 10
D30013 N30013 0 diode
R30014 N30013 N30014 10
D30014 N30014 0 diode
R30015 N30014 N30015 10
D30015 N30015 0 diode
R30016 N30015 N30016 10
D30016 N30016 0 diode
R30017 N30016 N30017 10
D30017 N30017 0 diode
R30018 N30017 N30018 10
D30018 N30018 0 diode
R30019 N30018 N30019 10
D30019 N30019 0 diode
R30020 N30019 N30020 10
D30020 N30020 0 diode
R30021 N30020 N30021 10
D30021 N30021 0 diode
R30022 N30021 N30022 10
D30022 N30022 0 diode
R30023 N30022 N30023 10
D30023 N30023 0 diode
R30024 N30023 N30024 10
D30024 N30024 0 diode
R30025 N30024 N30025 10
D30025 N30025 0 diode
R30026 N30025 N30026 10
D30026 N30026 0 diode
R30027 N30026 N30027 10
D30027 N30027 0 diode
R30028 N30027 N30028 10
D30028 N30028 0 diode
R30029 N30028 N30029 10
D30029 N30029 0 diode
R30030 N30029 N30030 10
D30030 N30030 0 diode
R30031 N30030 N30031 10
D30031 N30031 0 diode
R30032 N30031 N30032 10
D30032 N30032 0 diode
R30033 N30032 N30033 10
D30033 N30033 0 diode
R30034 N30033 N30034 10
D30034 N30034 0 diode
R30035 N30034 N30035 10
D30035 N30035 0 diode
R30036 N30035 N30036 10
D30036 N30036 0 diode
R30037 N30036 N30037 10
D30037 N30037 0 diode
R30038 N30037 N30038 10
D30038 N30038 0 diode
R30039 N30038 N30039 10
D30039 N30039 0 diode
R30040 N30039 N30040 10
D30040 N30040 0 diode
R30041 N30040 N30041 10
D30041 N30041 0 diode
R30042 N30041 N30042 10
D30042 N30042 0 diode
R30043 N30042 N30043 10
D30043 N30043 0 diode
R30044 N30043 N30044 10
D30044 N30044 0 diode
R30045 N30044 N30045 10
D30045 N30045 0 diode
R30046 N30045 N30046 10
D30046 N30046 0 diode
R30047 N30046 N30047 10
D30047 N30047 0 diode
R30048 N30047 N30048 10
D30048 N30048 0 diode
R30049 N30048 N30049 10
D30049 N30049 0 diode
R30050 N30049 N30050 10
D30050 N30050 0 diode
R30051 N30050 N30051 10
D30051 N30051 0 diode
R30052 N30051 N30052 10
D30052 N30052 0 diode
R30053 N30052 N30053 10
D30053 N30053 0 diode
R30054 N30053 N30054 10
D30054 N30054 0 diode
R30055 N30054 N30055 10
D30055 N30055 0 diode
R30056 N30055 N30056 10
D30056 N30056 0 diode
R30057 N30056 N30057 10
D30057 N30057 0 diode
R30058 N30057 N30058 10
D30058 N30058 0 diode
R30059 N30058 N30059 10
D30059 N30059 0 diode
R30060 N30059 N30060 10
D30060 N30060 0 diode
R30061 N30060 N30061 10
D30061 N30061 0 diode
R30062 N30061 N30062 10
D30062 N30062 0 diode
R30063 N30062 N30063 10
D30063 N30063 0 diode
R30064 N30063 N30064 10
D30064 N30064 0 diode
R30065 N30064 N30065 10
D30065 N30065 0 diode
R30066 N30065 N30066 10
D30066 N30066 0 diode
R30067 N30066 N30067 10
D30067 N30067 0 diode
R30068 N30067 N30068 10
D30068 N30068 0 diode
R30069 N30068 N30069 10
D30069 N30069 0 diode
R30070 N30069 N30070 10
D30070 N30070 0 diode
R30071 N30070 N30071 10
D30071 N30071 0 diode
R30072 N30071 N30072 10
D30072 N30072 0 diode
R30073 N30072 N30073 10
D30073 N30073 0 diode
R30074 N30073 N30074 10
D30074 N30074 0 diode
R30075 N30074 N30075 10
D30075 N30075 0 diode
R30076 N30075 N30076 10
D30076 N30076 0 diode
R30077 N30076 N30077 10
D30077 N30077 0 diode
R30078 N30077 N30078 10
D30078 N30078 0 diode
R30079 N30078 N30079 10
D30079 N30079 0 diode
R30080 N30079 N30080 10
D30080 N30080 0 diode
R30081 N30080 N30081 10
D30081 N30081 0 diode
R30082 N30081 N30082 10
D30082 N30082 0 diode
R30083 N30082 N30083 10
D30083 N30083 0 diode
R30084 N30083 N30084 10
D30084 N30084 0 diode
R30085 N30084 N30085 10
D30085 N30085 0 diode
R30086 N30085 N30086 10
D30086 N30086 0 diode
R30087 N30086 N30087 10
D30087 N30087 0 diode
R30088 N30087 N30088 10
D30088 N30088 0 diode
R30089 N30088 N30089 10
D30089 N30089 0 diode
R30090 N30089 N30090 10
D30090 N30090 0 diode
R30091 N30090 N30091 10
D30091 N30091 0 diode
R30092 N30091 N30092 10
D30092 N30092 0 diode
R30093 N30092 N30093 10
D30093 N30093 0 diode
R30094 N30093 N30094 10
D30094 N30094 0 diode
R30095 N30094 N30095 10
D30095 N30095 0 diode
R30096 N30095 N30096 10
D30096 N30096 0 diode
R30097 N30096 N30097 10
D30097 N30097 0 diode
R30098 N30097 N30098 10
D30098 N30098 0 diode
R30099 N30098 N30099 10
D30099 N30099 0 diode
R30100 N30099 N30100 10
D30100 N30100 0 diode
R30101 N30100 N30101 10
D30101 N30101 0 diode
R30102 N30101 N30102 10
D30102 N30102 0 diode
R30103 N30102 N30103 10
D30103 N30103 0 diode
R30104 N30103 N30104 10
D30104 N30104 0 diode
R30105 N30104 N30105 10
D30105 N30105 0 diode
R30106 N30105 N30106 10
D30106 N30106 0 diode
R30107 N30106 N30107 10
D30107 N30107 0 diode
R30108 N30107 N30108 10
D30108 N30108 0 diode
R30109 N30108 N30109 10
D30109 N30109 0 diode
R30110 N30109 N30110 10
D30110 N30110 0 diode
R30111 N30110 N30111 10
D30111 N30111 0 diode
R30112 N30111 N30112 10
D30112 N30112 0 diode
R30113 N30112 N30113 10
D30113 N30113 0 diode
R30114 N30113 N30114 10
D30114 N30114 0 diode
R30115 N30114 N30115 10
D30115 N30115 0 diode
R30116 N30115 N30116 10
D30116 N30116 0 diode
R30117 N30116 N30117 10
D30117 N30117 0 diode
R30118 N30117 N30118 10
D30118 N30118 0 diode
R30119 N30118 N30119 10
D30119 N30119 0 diode
R30120 N30119 N30120 10
D30120 N30120 0 diode
R30121 N30120 N30121 10
D30121 N30121 0 diode
R30122 N30121 N30122 10
D30122 N30122 0 diode
R30123 N30122 N30123 10
D30123 N30123 0 diode
R30124 N30123 N30124 10
D30124 N30124 0 diode
R30125 N30124 N30125 10
D30125 N30125 0 diode
R30126 N30125 N30126 10
D30126 N30126 0 diode
R30127 N30126 N30127 10
D30127 N30127 0 diode
R30128 N30127 N30128 10
D30128 N30128 0 diode
R30129 N30128 N30129 10
D30129 N30129 0 diode
R30130 N30129 N30130 10
D30130 N30130 0 diode
R30131 N30130 N30131 10
D30131 N30131 0 diode
R30132 N30131 N30132 10
D30132 N30132 0 diode
R30133 N30132 N30133 10
D30133 N30133 0 diode
R30134 N30133 N30134 10
D30134 N30134 0 diode
R30135 N30134 N30135 10
D30135 N30135 0 diode
R30136 N30135 N30136 10
D30136 N30136 0 diode
R30137 N30136 N30137 10
D30137 N30137 0 diode
R30138 N30137 N30138 10
D30138 N30138 0 diode
R30139 N30138 N30139 10
D30139 N30139 0 diode
R30140 N30139 N30140 10
D30140 N30140 0 diode
R30141 N30140 N30141 10
D30141 N30141 0 diode
R30142 N30141 N30142 10
D30142 N30142 0 diode
R30143 N30142 N30143 10
D30143 N30143 0 diode
R30144 N30143 N30144 10
D30144 N30144 0 diode
R30145 N30144 N30145 10
D30145 N30145 0 diode
R30146 N30145 N30146 10
D30146 N30146 0 diode
R30147 N30146 N30147 10
D30147 N30147 0 diode
R30148 N30147 N30148 10
D30148 N30148 0 diode
R30149 N30148 N30149 10
D30149 N30149 0 diode
R30150 N30149 N30150 10
D30150 N30150 0 diode
R30151 N30150 N30151 10
D30151 N30151 0 diode
R30152 N30151 N30152 10
D30152 N30152 0 diode
R30153 N30152 N30153 10
D30153 N30153 0 diode
R30154 N30153 N30154 10
D30154 N30154 0 diode
R30155 N30154 N30155 10
D30155 N30155 0 diode
R30156 N30155 N30156 10
D30156 N30156 0 diode
R30157 N30156 N30157 10
D30157 N30157 0 diode
R30158 N30157 N30158 10
D30158 N30158 0 diode
R30159 N30158 N30159 10
D30159 N30159 0 diode
R30160 N30159 N30160 10
D30160 N30160 0 diode
R30161 N30160 N30161 10
D30161 N30161 0 diode
R30162 N30161 N30162 10
D30162 N30162 0 diode
R30163 N30162 N30163 10
D30163 N30163 0 diode
R30164 N30163 N30164 10
D30164 N30164 0 diode
R30165 N30164 N30165 10
D30165 N30165 0 diode
R30166 N30165 N30166 10
D30166 N30166 0 diode
R30167 N30166 N30167 10
D30167 N30167 0 diode
R30168 N30167 N30168 10
D30168 N30168 0 diode
R30169 N30168 N30169 10
D30169 N30169 0 diode
R30170 N30169 N30170 10
D30170 N30170 0 diode
R30171 N30170 N30171 10
D30171 N30171 0 diode
R30172 N30171 N30172 10
D30172 N30172 0 diode
R30173 N30172 N30173 10
D30173 N30173 0 diode
R30174 N30173 N30174 10
D30174 N30174 0 diode
R30175 N30174 N30175 10
D30175 N30175 0 diode
R30176 N30175 N30176 10
D30176 N30176 0 diode
R30177 N30176 N30177 10
D30177 N30177 0 diode
R30178 N30177 N30178 10
D30178 N30178 0 diode
R30179 N30178 N30179 10
D30179 N30179 0 diode
R30180 N30179 N30180 10
D30180 N30180 0 diode
R30181 N30180 N30181 10
D30181 N30181 0 diode
R30182 N30181 N30182 10
D30182 N30182 0 diode
R30183 N30182 N30183 10
D30183 N30183 0 diode
R30184 N30183 N30184 10
D30184 N30184 0 diode
R30185 N30184 N30185 10
D30185 N30185 0 diode
R30186 N30185 N30186 10
D30186 N30186 0 diode
R30187 N30186 N30187 10
D30187 N30187 0 diode
R30188 N30187 N30188 10
D30188 N30188 0 diode
R30189 N30188 N30189 10
D30189 N30189 0 diode
R30190 N30189 N30190 10
D30190 N30190 0 diode
R30191 N30190 N30191 10
D30191 N30191 0 diode
R30192 N30191 N30192 10
D30192 N30192 0 diode
R30193 N30192 N30193 10
D30193 N30193 0 diode
R30194 N30193 N30194 10
D30194 N30194 0 diode
R30195 N30194 N30195 10
D30195 N30195 0 diode
R30196 N30195 N30196 10
D30196 N30196 0 diode
R30197 N30196 N30197 10
D30197 N30197 0 diode
R30198 N30197 N30198 10
D30198 N30198 0 diode
R30199 N30198 N30199 10
D30199 N30199 0 diode
R30200 N30199 N30200 10
D30200 N30200 0 diode
R30201 N30200 N30201 10
D30201 N30201 0 diode
R30202 N30201 N30202 10
D30202 N30202 0 diode
R30203 N30202 N30203 10
D30203 N30203 0 diode
R30204 N30203 N30204 10
D30204 N30204 0 diode
R30205 N30204 N30205 10
D30205 N30205 0 diode
R30206 N30205 N30206 10
D30206 N30206 0 diode
R30207 N30206 N30207 10
D30207 N30207 0 diode
R30208 N30207 N30208 10
D30208 N30208 0 diode
R30209 N30208 N30209 10
D30209 N30209 0 diode
R30210 N30209 N30210 10
D30210 N30210 0 diode
R30211 N30210 N30211 10
D30211 N30211 0 diode
R30212 N30211 N30212 10
D30212 N30212 0 diode
R30213 N30212 N30213 10
D30213 N30213 0 diode
R30214 N30213 N30214 10
D30214 N30214 0 diode
R30215 N30214 N30215 10
D30215 N30215 0 diode
R30216 N30215 N30216 10
D30216 N30216 0 diode
R30217 N30216 N30217 10
D30217 N30217 0 diode
R30218 N30217 N30218 10
D30218 N30218 0 diode
R30219 N30218 N30219 10
D30219 N30219 0 diode
R30220 N30219 N30220 10
D30220 N30220 0 diode
R30221 N30220 N30221 10
D30221 N30221 0 diode
R30222 N30221 N30222 10
D30222 N30222 0 diode
R30223 N30222 N30223 10
D30223 N30223 0 diode
R30224 N30223 N30224 10
D30224 N30224 0 diode
R30225 N30224 N30225 10
D30225 N30225 0 diode
R30226 N30225 N30226 10
D30226 N30226 0 diode
R30227 N30226 N30227 10
D30227 N30227 0 diode
R30228 N30227 N30228 10
D30228 N30228 0 diode
R30229 N30228 N30229 10
D30229 N30229 0 diode
R30230 N30229 N30230 10
D30230 N30230 0 diode
R30231 N30230 N30231 10
D30231 N30231 0 diode
R30232 N30231 N30232 10
D30232 N30232 0 diode
R30233 N30232 N30233 10
D30233 N30233 0 diode
R30234 N30233 N30234 10
D30234 N30234 0 diode
R30235 N30234 N30235 10
D30235 N30235 0 diode
R30236 N30235 N30236 10
D30236 N30236 0 diode
R30237 N30236 N30237 10
D30237 N30237 0 diode
R30238 N30237 N30238 10
D30238 N30238 0 diode
R30239 N30238 N30239 10
D30239 N30239 0 diode
R30240 N30239 N30240 10
D30240 N30240 0 diode
R30241 N30240 N30241 10
D30241 N30241 0 diode
R30242 N30241 N30242 10
D30242 N30242 0 diode
R30243 N30242 N30243 10
D30243 N30243 0 diode
R30244 N30243 N30244 10
D30244 N30244 0 diode
R30245 N30244 N30245 10
D30245 N30245 0 diode
R30246 N30245 N30246 10
D30246 N30246 0 diode
R30247 N30246 N30247 10
D30247 N30247 0 diode
R30248 N30247 N30248 10
D30248 N30248 0 diode
R30249 N30248 N30249 10
D30249 N30249 0 diode
R30250 N30249 N30250 10
D30250 N30250 0 diode
R30251 N30250 N30251 10
D30251 N30251 0 diode
R30252 N30251 N30252 10
D30252 N30252 0 diode
R30253 N30252 N30253 10
D30253 N30253 0 diode
R30254 N30253 N30254 10
D30254 N30254 0 diode
R30255 N30254 N30255 10
D30255 N30255 0 diode
R30256 N30255 N30256 10
D30256 N30256 0 diode
R30257 N30256 N30257 10
D30257 N30257 0 diode
R30258 N30257 N30258 10
D30258 N30258 0 diode
R30259 N30258 N30259 10
D30259 N30259 0 diode
R30260 N30259 N30260 10
D30260 N30260 0 diode
R30261 N30260 N30261 10
D30261 N30261 0 diode
R30262 N30261 N30262 10
D30262 N30262 0 diode
R30263 N30262 N30263 10
D30263 N30263 0 diode
R30264 N30263 N30264 10
D30264 N30264 0 diode
R30265 N30264 N30265 10
D30265 N30265 0 diode
R30266 N30265 N30266 10
D30266 N30266 0 diode
R30267 N30266 N30267 10
D30267 N30267 0 diode
R30268 N30267 N30268 10
D30268 N30268 0 diode
R30269 N30268 N30269 10
D30269 N30269 0 diode
R30270 N30269 N30270 10
D30270 N30270 0 diode
R30271 N30270 N30271 10
D30271 N30271 0 diode
R30272 N30271 N30272 10
D30272 N30272 0 diode
R30273 N30272 N30273 10
D30273 N30273 0 diode
R30274 N30273 N30274 10
D30274 N30274 0 diode
R30275 N30274 N30275 10
D30275 N30275 0 diode
R30276 N30275 N30276 10
D30276 N30276 0 diode
R30277 N30276 N30277 10
D30277 N30277 0 diode
R30278 N30277 N30278 10
D30278 N30278 0 diode
R30279 N30278 N30279 10
D30279 N30279 0 diode
R30280 N30279 N30280 10
D30280 N30280 0 diode
R30281 N30280 N30281 10
D30281 N30281 0 diode
R30282 N30281 N30282 10
D30282 N30282 0 diode
R30283 N30282 N30283 10
D30283 N30283 0 diode
R30284 N30283 N30284 10
D30284 N30284 0 diode
R30285 N30284 N30285 10
D30285 N30285 0 diode
R30286 N30285 N30286 10
D30286 N30286 0 diode
R30287 N30286 N30287 10
D30287 N30287 0 diode
R30288 N30287 N30288 10
D30288 N30288 0 diode
R30289 N30288 N30289 10
D30289 N30289 0 diode
R30290 N30289 N30290 10
D30290 N30290 0 diode
R30291 N30290 N30291 10
D30291 N30291 0 diode
R30292 N30291 N30292 10
D30292 N30292 0 diode
R30293 N30292 N30293 10
D30293 N30293 0 diode
R30294 N30293 N30294 10
D30294 N30294 0 diode
R30295 N30294 N30295 10
D30295 N30295 0 diode
R30296 N30295 N30296 10
D30296 N30296 0 diode
R30297 N30296 N30297 10
D30297 N30297 0 diode
R30298 N30297 N30298 10
D30298 N30298 0 diode
R30299 N30298 N30299 10
D30299 N30299 0 diode
R30300 N30299 N30300 10
D30300 N30300 0 diode
R30301 N30300 N30301 10
D30301 N30301 0 diode
R30302 N30301 N30302 10
D30302 N30302 0 diode
R30303 N30302 N30303 10
D30303 N30303 0 diode
R30304 N30303 N30304 10
D30304 N30304 0 diode
R30305 N30304 N30305 10
D30305 N30305 0 diode
R30306 N30305 N30306 10
D30306 N30306 0 diode
R30307 N30306 N30307 10
D30307 N30307 0 diode
R30308 N30307 N30308 10
D30308 N30308 0 diode
R30309 N30308 N30309 10
D30309 N30309 0 diode
R30310 N30309 N30310 10
D30310 N30310 0 diode
R30311 N30310 N30311 10
D30311 N30311 0 diode
R30312 N30311 N30312 10
D30312 N30312 0 diode
R30313 N30312 N30313 10
D30313 N30313 0 diode
R30314 N30313 N30314 10
D30314 N30314 0 diode
R30315 N30314 N30315 10
D30315 N30315 0 diode
R30316 N30315 N30316 10
D30316 N30316 0 diode
R30317 N30316 N30317 10
D30317 N30317 0 diode
R30318 N30317 N30318 10
D30318 N30318 0 diode
R30319 N30318 N30319 10
D30319 N30319 0 diode
R30320 N30319 N30320 10
D30320 N30320 0 diode
R30321 N30320 N30321 10
D30321 N30321 0 diode
R30322 N30321 N30322 10
D30322 N30322 0 diode
R30323 N30322 N30323 10
D30323 N30323 0 diode
R30324 N30323 N30324 10
D30324 N30324 0 diode
R30325 N30324 N30325 10
D30325 N30325 0 diode
R30326 N30325 N30326 10
D30326 N30326 0 diode
R30327 N30326 N30327 10
D30327 N30327 0 diode
R30328 N30327 N30328 10
D30328 N30328 0 diode
R30329 N30328 N30329 10
D30329 N30329 0 diode
R30330 N30329 N30330 10
D30330 N30330 0 diode
R30331 N30330 N30331 10
D30331 N30331 0 diode
R30332 N30331 N30332 10
D30332 N30332 0 diode
R30333 N30332 N30333 10
D30333 N30333 0 diode
R30334 N30333 N30334 10
D30334 N30334 0 diode
R30335 N30334 N30335 10
D30335 N30335 0 diode
R30336 N30335 N30336 10
D30336 N30336 0 diode
R30337 N30336 N30337 10
D30337 N30337 0 diode
R30338 N30337 N30338 10
D30338 N30338 0 diode
R30339 N30338 N30339 10
D30339 N30339 0 diode
R30340 N30339 N30340 10
D30340 N30340 0 diode
R30341 N30340 N30341 10
D30341 N30341 0 diode
R30342 N30341 N30342 10
D30342 N30342 0 diode
R30343 N30342 N30343 10
D30343 N30343 0 diode
R30344 N30343 N30344 10
D30344 N30344 0 diode
R30345 N30344 N30345 10
D30345 N30345 0 diode
R30346 N30345 N30346 10
D30346 N30346 0 diode
R30347 N30346 N30347 10
D30347 N30347 0 diode
R30348 N30347 N30348 10
D30348 N30348 0 diode
R30349 N30348 N30349 10
D30349 N30349 0 diode
R30350 N30349 N30350 10
D30350 N30350 0 diode
R30351 N30350 N30351 10
D30351 N30351 0 diode
R30352 N30351 N30352 10
D30352 N30352 0 diode
R30353 N30352 N30353 10
D30353 N30353 0 diode
R30354 N30353 N30354 10
D30354 N30354 0 diode
R30355 N30354 N30355 10
D30355 N30355 0 diode
R30356 N30355 N30356 10
D30356 N30356 0 diode
R30357 N30356 N30357 10
D30357 N30357 0 diode
R30358 N30357 N30358 10
D30358 N30358 0 diode
R30359 N30358 N30359 10
D30359 N30359 0 diode
R30360 N30359 N30360 10
D30360 N30360 0 diode
R30361 N30360 N30361 10
D30361 N30361 0 diode
R30362 N30361 N30362 10
D30362 N30362 0 diode
R30363 N30362 N30363 10
D30363 N30363 0 diode
R30364 N30363 N30364 10
D30364 N30364 0 diode
R30365 N30364 N30365 10
D30365 N30365 0 diode
R30366 N30365 N30366 10
D30366 N30366 0 diode
R30367 N30366 N30367 10
D30367 N30367 0 diode
R30368 N30367 N30368 10
D30368 N30368 0 diode
R30369 N30368 N30369 10
D30369 N30369 0 diode
R30370 N30369 N30370 10
D30370 N30370 0 diode
R30371 N30370 N30371 10
D30371 N30371 0 diode
R30372 N30371 N30372 10
D30372 N30372 0 diode
R30373 N30372 N30373 10
D30373 N30373 0 diode
R30374 N30373 N30374 10
D30374 N30374 0 diode
R30375 N30374 N30375 10
D30375 N30375 0 diode
R30376 N30375 N30376 10
D30376 N30376 0 diode
R30377 N30376 N30377 10
D30377 N30377 0 diode
R30378 N30377 N30378 10
D30378 N30378 0 diode
R30379 N30378 N30379 10
D30379 N30379 0 diode
R30380 N30379 N30380 10
D30380 N30380 0 diode
R30381 N30380 N30381 10
D30381 N30381 0 diode
R30382 N30381 N30382 10
D30382 N30382 0 diode
R30383 N30382 N30383 10
D30383 N30383 0 diode
R30384 N30383 N30384 10
D30384 N30384 0 diode
R30385 N30384 N30385 10
D30385 N30385 0 diode
R30386 N30385 N30386 10
D30386 N30386 0 diode
R30387 N30386 N30387 10
D30387 N30387 0 diode
R30388 N30387 N30388 10
D30388 N30388 0 diode
R30389 N30388 N30389 10
D30389 N30389 0 diode
R30390 N30389 N30390 10
D30390 N30390 0 diode
R30391 N30390 N30391 10
D30391 N30391 0 diode
R30392 N30391 N30392 10
D30392 N30392 0 diode
R30393 N30392 N30393 10
D30393 N30393 0 diode
R30394 N30393 N30394 10
D30394 N30394 0 diode
R30395 N30394 N30395 10
D30395 N30395 0 diode
R30396 N30395 N30396 10
D30396 N30396 0 diode
R30397 N30396 N30397 10
D30397 N30397 0 diode
R30398 N30397 N30398 10
D30398 N30398 0 diode
R30399 N30398 N30399 10
D30399 N30399 0 diode
R30400 N30399 N30400 10
D30400 N30400 0 diode
R30401 N30400 N30401 10
D30401 N30401 0 diode
R30402 N30401 N30402 10
D30402 N30402 0 diode
R30403 N30402 N30403 10
D30403 N30403 0 diode
R30404 N30403 N30404 10
D30404 N30404 0 diode
R30405 N30404 N30405 10
D30405 N30405 0 diode
R30406 N30405 N30406 10
D30406 N30406 0 diode
R30407 N30406 N30407 10
D30407 N30407 0 diode
R30408 N30407 N30408 10
D30408 N30408 0 diode
R30409 N30408 N30409 10
D30409 N30409 0 diode
R30410 N30409 N30410 10
D30410 N30410 0 diode
R30411 N30410 N30411 10
D30411 N30411 0 diode
R30412 N30411 N30412 10
D30412 N30412 0 diode
R30413 N30412 N30413 10
D30413 N30413 0 diode
R30414 N30413 N30414 10
D30414 N30414 0 diode
R30415 N30414 N30415 10
D30415 N30415 0 diode
R30416 N30415 N30416 10
D30416 N30416 0 diode
R30417 N30416 N30417 10
D30417 N30417 0 diode
R30418 N30417 N30418 10
D30418 N30418 0 diode
R30419 N30418 N30419 10
D30419 N30419 0 diode
R30420 N30419 N30420 10
D30420 N30420 0 diode
R30421 N30420 N30421 10
D30421 N30421 0 diode
R30422 N30421 N30422 10
D30422 N30422 0 diode
R30423 N30422 N30423 10
D30423 N30423 0 diode
R30424 N30423 N30424 10
D30424 N30424 0 diode
R30425 N30424 N30425 10
D30425 N30425 0 diode
R30426 N30425 N30426 10
D30426 N30426 0 diode
R30427 N30426 N30427 10
D30427 N30427 0 diode
R30428 N30427 N30428 10
D30428 N30428 0 diode
R30429 N30428 N30429 10
D30429 N30429 0 diode
R30430 N30429 N30430 10
D30430 N30430 0 diode
R30431 N30430 N30431 10
D30431 N30431 0 diode
R30432 N30431 N30432 10
D30432 N30432 0 diode
R30433 N30432 N30433 10
D30433 N30433 0 diode
R30434 N30433 N30434 10
D30434 N30434 0 diode
R30435 N30434 N30435 10
D30435 N30435 0 diode
R30436 N30435 N30436 10
D30436 N30436 0 diode
R30437 N30436 N30437 10
D30437 N30437 0 diode
R30438 N30437 N30438 10
D30438 N30438 0 diode
R30439 N30438 N30439 10
D30439 N30439 0 diode
R30440 N30439 N30440 10
D30440 N30440 0 diode
R30441 N30440 N30441 10
D30441 N30441 0 diode
R30442 N30441 N30442 10
D30442 N30442 0 diode
R30443 N30442 N30443 10
D30443 N30443 0 diode
R30444 N30443 N30444 10
D30444 N30444 0 diode
R30445 N30444 N30445 10
D30445 N30445 0 diode
R30446 N30445 N30446 10
D30446 N30446 0 diode
R30447 N30446 N30447 10
D30447 N30447 0 diode
R30448 N30447 N30448 10
D30448 N30448 0 diode
R30449 N30448 N30449 10
D30449 N30449 0 diode
R30450 N30449 N30450 10
D30450 N30450 0 diode
R30451 N30450 N30451 10
D30451 N30451 0 diode
R30452 N30451 N30452 10
D30452 N30452 0 diode
R30453 N30452 N30453 10
D30453 N30453 0 diode
R30454 N30453 N30454 10
D30454 N30454 0 diode
R30455 N30454 N30455 10
D30455 N30455 0 diode
R30456 N30455 N30456 10
D30456 N30456 0 diode
R30457 N30456 N30457 10
D30457 N30457 0 diode
R30458 N30457 N30458 10
D30458 N30458 0 diode
R30459 N30458 N30459 10
D30459 N30459 0 diode
R30460 N30459 N30460 10
D30460 N30460 0 diode
R30461 N30460 N30461 10
D30461 N30461 0 diode
R30462 N30461 N30462 10
D30462 N30462 0 diode
R30463 N30462 N30463 10
D30463 N30463 0 diode
R30464 N30463 N30464 10
D30464 N30464 0 diode
R30465 N30464 N30465 10
D30465 N30465 0 diode
R30466 N30465 N30466 10
D30466 N30466 0 diode
R30467 N30466 N30467 10
D30467 N30467 0 diode
R30468 N30467 N30468 10
D30468 N30468 0 diode
R30469 N30468 N30469 10
D30469 N30469 0 diode
R30470 N30469 N30470 10
D30470 N30470 0 diode
R30471 N30470 N30471 10
D30471 N30471 0 diode
R30472 N30471 N30472 10
D30472 N30472 0 diode
R30473 N30472 N30473 10
D30473 N30473 0 diode
R30474 N30473 N30474 10
D30474 N30474 0 diode
R30475 N30474 N30475 10
D30475 N30475 0 diode
R30476 N30475 N30476 10
D30476 N30476 0 diode
R30477 N30476 N30477 10
D30477 N30477 0 diode
R30478 N30477 N30478 10
D30478 N30478 0 diode
R30479 N30478 N30479 10
D30479 N30479 0 diode
R30480 N30479 N30480 10
D30480 N30480 0 diode
R30481 N30480 N30481 10
D30481 N30481 0 diode
R30482 N30481 N30482 10
D30482 N30482 0 diode
R30483 N30482 N30483 10
D30483 N30483 0 diode
R30484 N30483 N30484 10
D30484 N30484 0 diode
R30485 N30484 N30485 10
D30485 N30485 0 diode
R30486 N30485 N30486 10
D30486 N30486 0 diode
R30487 N30486 N30487 10
D30487 N30487 0 diode
R30488 N30487 N30488 10
D30488 N30488 0 diode
R30489 N30488 N30489 10
D30489 N30489 0 diode
R30490 N30489 N30490 10
D30490 N30490 0 diode
R30491 N30490 N30491 10
D30491 N30491 0 diode
R30492 N30491 N30492 10
D30492 N30492 0 diode
R30493 N30492 N30493 10
D30493 N30493 0 diode
R30494 N30493 N30494 10
D30494 N30494 0 diode
R30495 N30494 N30495 10
D30495 N30495 0 diode
R30496 N30495 N30496 10
D30496 N30496 0 diode
R30497 N30496 N30497 10
D30497 N30497 0 diode
R30498 N30497 N30498 10
D30498 N30498 0 diode
R30499 N30498 N30499 10
D30499 N30499 0 diode
R30500 N30499 N30500 10
D30500 N30500 0 diode
R30501 N30500 N30501 10
D30501 N30501 0 diode
R30502 N30501 N30502 10
D30502 N30502 0 diode
R30503 N30502 N30503 10
D30503 N30503 0 diode
R30504 N30503 N30504 10
D30504 N30504 0 diode
R30505 N30504 N30505 10
D30505 N30505 0 diode
R30506 N30505 N30506 10
D30506 N30506 0 diode
R30507 N30506 N30507 10
D30507 N30507 0 diode
R30508 N30507 N30508 10
D30508 N30508 0 diode
R30509 N30508 N30509 10
D30509 N30509 0 diode
R30510 N30509 N30510 10
D30510 N30510 0 diode
R30511 N30510 N30511 10
D30511 N30511 0 diode
R30512 N30511 N30512 10
D30512 N30512 0 diode
R30513 N30512 N30513 10
D30513 N30513 0 diode
R30514 N30513 N30514 10
D30514 N30514 0 diode
R30515 N30514 N30515 10
D30515 N30515 0 diode
R30516 N30515 N30516 10
D30516 N30516 0 diode
R30517 N30516 N30517 10
D30517 N30517 0 diode
R30518 N30517 N30518 10
D30518 N30518 0 diode
R30519 N30518 N30519 10
D30519 N30519 0 diode
R30520 N30519 N30520 10
D30520 N30520 0 diode
R30521 N30520 N30521 10
D30521 N30521 0 diode
R30522 N30521 N30522 10
D30522 N30522 0 diode
R30523 N30522 N30523 10
D30523 N30523 0 diode
R30524 N30523 N30524 10
D30524 N30524 0 diode
R30525 N30524 N30525 10
D30525 N30525 0 diode
R30526 N30525 N30526 10
D30526 N30526 0 diode
R30527 N30526 N30527 10
D30527 N30527 0 diode
R30528 N30527 N30528 10
D30528 N30528 0 diode
R30529 N30528 N30529 10
D30529 N30529 0 diode
R30530 N30529 N30530 10
D30530 N30530 0 diode
R30531 N30530 N30531 10
D30531 N30531 0 diode
R30532 N30531 N30532 10
D30532 N30532 0 diode
R30533 N30532 N30533 10
D30533 N30533 0 diode
R30534 N30533 N30534 10
D30534 N30534 0 diode
R30535 N30534 N30535 10
D30535 N30535 0 diode
R30536 N30535 N30536 10
D30536 N30536 0 diode
R30537 N30536 N30537 10
D30537 N30537 0 diode
R30538 N30537 N30538 10
D30538 N30538 0 diode
R30539 N30538 N30539 10
D30539 N30539 0 diode
R30540 N30539 N30540 10
D30540 N30540 0 diode
R30541 N30540 N30541 10
D30541 N30541 0 diode
R30542 N30541 N30542 10
D30542 N30542 0 diode
R30543 N30542 N30543 10
D30543 N30543 0 diode
R30544 N30543 N30544 10
D30544 N30544 0 diode
R30545 N30544 N30545 10
D30545 N30545 0 diode
R30546 N30545 N30546 10
D30546 N30546 0 diode
R30547 N30546 N30547 10
D30547 N30547 0 diode
R30548 N30547 N30548 10
D30548 N30548 0 diode
R30549 N30548 N30549 10
D30549 N30549 0 diode
R30550 N30549 N30550 10
D30550 N30550 0 diode
R30551 N30550 N30551 10
D30551 N30551 0 diode
R30552 N30551 N30552 10
D30552 N30552 0 diode
R30553 N30552 N30553 10
D30553 N30553 0 diode
R30554 N30553 N30554 10
D30554 N30554 0 diode
R30555 N30554 N30555 10
D30555 N30555 0 diode
R30556 N30555 N30556 10
D30556 N30556 0 diode
R30557 N30556 N30557 10
D30557 N30557 0 diode
R30558 N30557 N30558 10
D30558 N30558 0 diode
R30559 N30558 N30559 10
D30559 N30559 0 diode
R30560 N30559 N30560 10
D30560 N30560 0 diode
R30561 N30560 N30561 10
D30561 N30561 0 diode
R30562 N30561 N30562 10
D30562 N30562 0 diode
R30563 N30562 N30563 10
D30563 N30563 0 diode
R30564 N30563 N30564 10
D30564 N30564 0 diode
R30565 N30564 N30565 10
D30565 N30565 0 diode
R30566 N30565 N30566 10
D30566 N30566 0 diode
R30567 N30566 N30567 10
D30567 N30567 0 diode
R30568 N30567 N30568 10
D30568 N30568 0 diode
R30569 N30568 N30569 10
D30569 N30569 0 diode
R30570 N30569 N30570 10
D30570 N30570 0 diode
R30571 N30570 N30571 10
D30571 N30571 0 diode
R30572 N30571 N30572 10
D30572 N30572 0 diode
R30573 N30572 N30573 10
D30573 N30573 0 diode
R30574 N30573 N30574 10
D30574 N30574 0 diode
R30575 N30574 N30575 10
D30575 N30575 0 diode
R30576 N30575 N30576 10
D30576 N30576 0 diode
R30577 N30576 N30577 10
D30577 N30577 0 diode
R30578 N30577 N30578 10
D30578 N30578 0 diode
R30579 N30578 N30579 10
D30579 N30579 0 diode
R30580 N30579 N30580 10
D30580 N30580 0 diode
R30581 N30580 N30581 10
D30581 N30581 0 diode
R30582 N30581 N30582 10
D30582 N30582 0 diode
R30583 N30582 N30583 10
D30583 N30583 0 diode
R30584 N30583 N30584 10
D30584 N30584 0 diode
R30585 N30584 N30585 10
D30585 N30585 0 diode
R30586 N30585 N30586 10
D30586 N30586 0 diode
R30587 N30586 N30587 10
D30587 N30587 0 diode
R30588 N30587 N30588 10
D30588 N30588 0 diode
R30589 N30588 N30589 10
D30589 N30589 0 diode
R30590 N30589 N30590 10
D30590 N30590 0 diode
R30591 N30590 N30591 10
D30591 N30591 0 diode
R30592 N30591 N30592 10
D30592 N30592 0 diode
R30593 N30592 N30593 10
D30593 N30593 0 diode
R30594 N30593 N30594 10
D30594 N30594 0 diode
R30595 N30594 N30595 10
D30595 N30595 0 diode
R30596 N30595 N30596 10
D30596 N30596 0 diode
R30597 N30596 N30597 10
D30597 N30597 0 diode
R30598 N30597 N30598 10
D30598 N30598 0 diode
R30599 N30598 N30599 10
D30599 N30599 0 diode
R30600 N30599 N30600 10
D30600 N30600 0 diode
R30601 N30600 N30601 10
D30601 N30601 0 diode
R30602 N30601 N30602 10
D30602 N30602 0 diode
R30603 N30602 N30603 10
D30603 N30603 0 diode
R30604 N30603 N30604 10
D30604 N30604 0 diode
R30605 N30604 N30605 10
D30605 N30605 0 diode
R30606 N30605 N30606 10
D30606 N30606 0 diode
R30607 N30606 N30607 10
D30607 N30607 0 diode
R30608 N30607 N30608 10
D30608 N30608 0 diode
R30609 N30608 N30609 10
D30609 N30609 0 diode
R30610 N30609 N30610 10
D30610 N30610 0 diode
R30611 N30610 N30611 10
D30611 N30611 0 diode
R30612 N30611 N30612 10
D30612 N30612 0 diode
R30613 N30612 N30613 10
D30613 N30613 0 diode
R30614 N30613 N30614 10
D30614 N30614 0 diode
R30615 N30614 N30615 10
D30615 N30615 0 diode
R30616 N30615 N30616 10
D30616 N30616 0 diode
R30617 N30616 N30617 10
D30617 N30617 0 diode
R30618 N30617 N30618 10
D30618 N30618 0 diode
R30619 N30618 N30619 10
D30619 N30619 0 diode
R30620 N30619 N30620 10
D30620 N30620 0 diode
R30621 N30620 N30621 10
D30621 N30621 0 diode
R30622 N30621 N30622 10
D30622 N30622 0 diode
R30623 N30622 N30623 10
D30623 N30623 0 diode
R30624 N30623 N30624 10
D30624 N30624 0 diode
R30625 N30624 N30625 10
D30625 N30625 0 diode
R30626 N30625 N30626 10
D30626 N30626 0 diode
R30627 N30626 N30627 10
D30627 N30627 0 diode
R30628 N30627 N30628 10
D30628 N30628 0 diode
R30629 N30628 N30629 10
D30629 N30629 0 diode
R30630 N30629 N30630 10
D30630 N30630 0 diode
R30631 N30630 N30631 10
D30631 N30631 0 diode
R30632 N30631 N30632 10
D30632 N30632 0 diode
R30633 N30632 N30633 10
D30633 N30633 0 diode
R30634 N30633 N30634 10
D30634 N30634 0 diode
R30635 N30634 N30635 10
D30635 N30635 0 diode
R30636 N30635 N30636 10
D30636 N30636 0 diode
R30637 N30636 N30637 10
D30637 N30637 0 diode
R30638 N30637 N30638 10
D30638 N30638 0 diode
R30639 N30638 N30639 10
D30639 N30639 0 diode
R30640 N30639 N30640 10
D30640 N30640 0 diode
R30641 N30640 N30641 10
D30641 N30641 0 diode
R30642 N30641 N30642 10
D30642 N30642 0 diode
R30643 N30642 N30643 10
D30643 N30643 0 diode
R30644 N30643 N30644 10
D30644 N30644 0 diode
R30645 N30644 N30645 10
D30645 N30645 0 diode
R30646 N30645 N30646 10
D30646 N30646 0 diode
R30647 N30646 N30647 10
D30647 N30647 0 diode
R30648 N30647 N30648 10
D30648 N30648 0 diode
R30649 N30648 N30649 10
D30649 N30649 0 diode
R30650 N30649 N30650 10
D30650 N30650 0 diode
R30651 N30650 N30651 10
D30651 N30651 0 diode
R30652 N30651 N30652 10
D30652 N30652 0 diode
R30653 N30652 N30653 10
D30653 N30653 0 diode
R30654 N30653 N30654 10
D30654 N30654 0 diode
R30655 N30654 N30655 10
D30655 N30655 0 diode
R30656 N30655 N30656 10
D30656 N30656 0 diode
R30657 N30656 N30657 10
D30657 N30657 0 diode
R30658 N30657 N30658 10
D30658 N30658 0 diode
R30659 N30658 N30659 10
D30659 N30659 0 diode
R30660 N30659 N30660 10
D30660 N30660 0 diode
R30661 N30660 N30661 10
D30661 N30661 0 diode
R30662 N30661 N30662 10
D30662 N30662 0 diode
R30663 N30662 N30663 10
D30663 N30663 0 diode
R30664 N30663 N30664 10
D30664 N30664 0 diode
R30665 N30664 N30665 10
D30665 N30665 0 diode
R30666 N30665 N30666 10
D30666 N30666 0 diode
R30667 N30666 N30667 10
D30667 N30667 0 diode
R30668 N30667 N30668 10
D30668 N30668 0 diode
R30669 N30668 N30669 10
D30669 N30669 0 diode
R30670 N30669 N30670 10
D30670 N30670 0 diode
R30671 N30670 N30671 10
D30671 N30671 0 diode
R30672 N30671 N30672 10
D30672 N30672 0 diode
R30673 N30672 N30673 10
D30673 N30673 0 diode
R30674 N30673 N30674 10
D30674 N30674 0 diode
R30675 N30674 N30675 10
D30675 N30675 0 diode
R30676 N30675 N30676 10
D30676 N30676 0 diode
R30677 N30676 N30677 10
D30677 N30677 0 diode
R30678 N30677 N30678 10
D30678 N30678 0 diode
R30679 N30678 N30679 10
D30679 N30679 0 diode
R30680 N30679 N30680 10
D30680 N30680 0 diode
R30681 N30680 N30681 10
D30681 N30681 0 diode
R30682 N30681 N30682 10
D30682 N30682 0 diode
R30683 N30682 N30683 10
D30683 N30683 0 diode
R30684 N30683 N30684 10
D30684 N30684 0 diode
R30685 N30684 N30685 10
D30685 N30685 0 diode
R30686 N30685 N30686 10
D30686 N30686 0 diode
R30687 N30686 N30687 10
D30687 N30687 0 diode
R30688 N30687 N30688 10
D30688 N30688 0 diode
R30689 N30688 N30689 10
D30689 N30689 0 diode
R30690 N30689 N30690 10
D30690 N30690 0 diode
R30691 N30690 N30691 10
D30691 N30691 0 diode
R30692 N30691 N30692 10
D30692 N30692 0 diode
R30693 N30692 N30693 10
D30693 N30693 0 diode
R30694 N30693 N30694 10
D30694 N30694 0 diode
R30695 N30694 N30695 10
D30695 N30695 0 diode
R30696 N30695 N30696 10
D30696 N30696 0 diode
R30697 N30696 N30697 10
D30697 N30697 0 diode
R30698 N30697 N30698 10
D30698 N30698 0 diode
R30699 N30698 N30699 10
D30699 N30699 0 diode
R30700 N30699 N30700 10
D30700 N30700 0 diode
R30701 N30700 N30701 10
D30701 N30701 0 diode
R30702 N30701 N30702 10
D30702 N30702 0 diode
R30703 N30702 N30703 10
D30703 N30703 0 diode
R30704 N30703 N30704 10
D30704 N30704 0 diode
R30705 N30704 N30705 10
D30705 N30705 0 diode
R30706 N30705 N30706 10
D30706 N30706 0 diode
R30707 N30706 N30707 10
D30707 N30707 0 diode
R30708 N30707 N30708 10
D30708 N30708 0 diode
R30709 N30708 N30709 10
D30709 N30709 0 diode
R30710 N30709 N30710 10
D30710 N30710 0 diode
R30711 N30710 N30711 10
D30711 N30711 0 diode
R30712 N30711 N30712 10
D30712 N30712 0 diode
R30713 N30712 N30713 10
D30713 N30713 0 diode
R30714 N30713 N30714 10
D30714 N30714 0 diode
R30715 N30714 N30715 10
D30715 N30715 0 diode
R30716 N30715 N30716 10
D30716 N30716 0 diode
R30717 N30716 N30717 10
D30717 N30717 0 diode
R30718 N30717 N30718 10
D30718 N30718 0 diode
R30719 N30718 N30719 10
D30719 N30719 0 diode
R30720 N30719 N30720 10
D30720 N30720 0 diode
R30721 N30720 N30721 10
D30721 N30721 0 diode
R30722 N30721 N30722 10
D30722 N30722 0 diode
R30723 N30722 N30723 10
D30723 N30723 0 diode
R30724 N30723 N30724 10
D30724 N30724 0 diode
R30725 N30724 N30725 10
D30725 N30725 0 diode
R30726 N30725 N30726 10
D30726 N30726 0 diode
R30727 N30726 N30727 10
D30727 N30727 0 diode
R30728 N30727 N30728 10
D30728 N30728 0 diode
R30729 N30728 N30729 10
D30729 N30729 0 diode
R30730 N30729 N30730 10
D30730 N30730 0 diode
R30731 N30730 N30731 10
D30731 N30731 0 diode
R30732 N30731 N30732 10
D30732 N30732 0 diode
R30733 N30732 N30733 10
D30733 N30733 0 diode
R30734 N30733 N30734 10
D30734 N30734 0 diode
R30735 N30734 N30735 10
D30735 N30735 0 diode
R30736 N30735 N30736 10
D30736 N30736 0 diode
R30737 N30736 N30737 10
D30737 N30737 0 diode
R30738 N30737 N30738 10
D30738 N30738 0 diode
R30739 N30738 N30739 10
D30739 N30739 0 diode
R30740 N30739 N30740 10
D30740 N30740 0 diode
R30741 N30740 N30741 10
D30741 N30741 0 diode
R30742 N30741 N30742 10
D30742 N30742 0 diode
R30743 N30742 N30743 10
D30743 N30743 0 diode
R30744 N30743 N30744 10
D30744 N30744 0 diode
R30745 N30744 N30745 10
D30745 N30745 0 diode
R30746 N30745 N30746 10
D30746 N30746 0 diode
R30747 N30746 N30747 10
D30747 N30747 0 diode
R30748 N30747 N30748 10
D30748 N30748 0 diode
R30749 N30748 N30749 10
D30749 N30749 0 diode
R30750 N30749 N30750 10
D30750 N30750 0 diode
R30751 N30750 N30751 10
D30751 N30751 0 diode
R30752 N30751 N30752 10
D30752 N30752 0 diode
R30753 N30752 N30753 10
D30753 N30753 0 diode
R30754 N30753 N30754 10
D30754 N30754 0 diode
R30755 N30754 N30755 10
D30755 N30755 0 diode
R30756 N30755 N30756 10
D30756 N30756 0 diode
R30757 N30756 N30757 10
D30757 N30757 0 diode
R30758 N30757 N30758 10
D30758 N30758 0 diode
R30759 N30758 N30759 10
D30759 N30759 0 diode
R30760 N30759 N30760 10
D30760 N30760 0 diode
R30761 N30760 N30761 10
D30761 N30761 0 diode
R30762 N30761 N30762 10
D30762 N30762 0 diode
R30763 N30762 N30763 10
D30763 N30763 0 diode
R30764 N30763 N30764 10
D30764 N30764 0 diode
R30765 N30764 N30765 10
D30765 N30765 0 diode
R30766 N30765 N30766 10
D30766 N30766 0 diode
R30767 N30766 N30767 10
D30767 N30767 0 diode
R30768 N30767 N30768 10
D30768 N30768 0 diode
R30769 N30768 N30769 10
D30769 N30769 0 diode
R30770 N30769 N30770 10
D30770 N30770 0 diode
R30771 N30770 N30771 10
D30771 N30771 0 diode
R30772 N30771 N30772 10
D30772 N30772 0 diode
R30773 N30772 N30773 10
D30773 N30773 0 diode
R30774 N30773 N30774 10
D30774 N30774 0 diode
R30775 N30774 N30775 10
D30775 N30775 0 diode
R30776 N30775 N30776 10
D30776 N30776 0 diode
R30777 N30776 N30777 10
D30777 N30777 0 diode
R30778 N30777 N30778 10
D30778 N30778 0 diode
R30779 N30778 N30779 10
D30779 N30779 0 diode
R30780 N30779 N30780 10
D30780 N30780 0 diode
R30781 N30780 N30781 10
D30781 N30781 0 diode
R30782 N30781 N30782 10
D30782 N30782 0 diode
R30783 N30782 N30783 10
D30783 N30783 0 diode
R30784 N30783 N30784 10
D30784 N30784 0 diode
R30785 N30784 N30785 10
D30785 N30785 0 diode
R30786 N30785 N30786 10
D30786 N30786 0 diode
R30787 N30786 N30787 10
D30787 N30787 0 diode
R30788 N30787 N30788 10
D30788 N30788 0 diode
R30789 N30788 N30789 10
D30789 N30789 0 diode
R30790 N30789 N30790 10
D30790 N30790 0 diode
R30791 N30790 N30791 10
D30791 N30791 0 diode
R30792 N30791 N30792 10
D30792 N30792 0 diode
R30793 N30792 N30793 10
D30793 N30793 0 diode
R30794 N30793 N30794 10
D30794 N30794 0 diode
R30795 N30794 N30795 10
D30795 N30795 0 diode
R30796 N30795 N30796 10
D30796 N30796 0 diode
R30797 N30796 N30797 10
D30797 N30797 0 diode
R30798 N30797 N30798 10
D30798 N30798 0 diode
R30799 N30798 N30799 10
D30799 N30799 0 diode
R30800 N30799 N30800 10
D30800 N30800 0 diode
R30801 N30800 N30801 10
D30801 N30801 0 diode
R30802 N30801 N30802 10
D30802 N30802 0 diode
R30803 N30802 N30803 10
D30803 N30803 0 diode
R30804 N30803 N30804 10
D30804 N30804 0 diode
R30805 N30804 N30805 10
D30805 N30805 0 diode
R30806 N30805 N30806 10
D30806 N30806 0 diode
R30807 N30806 N30807 10
D30807 N30807 0 diode
R30808 N30807 N30808 10
D30808 N30808 0 diode
R30809 N30808 N30809 10
D30809 N30809 0 diode
R30810 N30809 N30810 10
D30810 N30810 0 diode
R30811 N30810 N30811 10
D30811 N30811 0 diode
R30812 N30811 N30812 10
D30812 N30812 0 diode
R30813 N30812 N30813 10
D30813 N30813 0 diode
R30814 N30813 N30814 10
D30814 N30814 0 diode
R30815 N30814 N30815 10
D30815 N30815 0 diode
R30816 N30815 N30816 10
D30816 N30816 0 diode
R30817 N30816 N30817 10
D30817 N30817 0 diode
R30818 N30817 N30818 10
D30818 N30818 0 diode
R30819 N30818 N30819 10
D30819 N30819 0 diode
R30820 N30819 N30820 10
D30820 N30820 0 diode
R30821 N30820 N30821 10
D30821 N30821 0 diode
R30822 N30821 N30822 10
D30822 N30822 0 diode
R30823 N30822 N30823 10
D30823 N30823 0 diode
R30824 N30823 N30824 10
D30824 N30824 0 diode
R30825 N30824 N30825 10
D30825 N30825 0 diode
R30826 N30825 N30826 10
D30826 N30826 0 diode
R30827 N30826 N30827 10
D30827 N30827 0 diode
R30828 N30827 N30828 10
D30828 N30828 0 diode
R30829 N30828 N30829 10
D30829 N30829 0 diode
R30830 N30829 N30830 10
D30830 N30830 0 diode
R30831 N30830 N30831 10
D30831 N30831 0 diode
R30832 N30831 N30832 10
D30832 N30832 0 diode
R30833 N30832 N30833 10
D30833 N30833 0 diode
R30834 N30833 N30834 10
D30834 N30834 0 diode
R30835 N30834 N30835 10
D30835 N30835 0 diode
R30836 N30835 N30836 10
D30836 N30836 0 diode
R30837 N30836 N30837 10
D30837 N30837 0 diode
R30838 N30837 N30838 10
D30838 N30838 0 diode
R30839 N30838 N30839 10
D30839 N30839 0 diode
R30840 N30839 N30840 10
D30840 N30840 0 diode
R30841 N30840 N30841 10
D30841 N30841 0 diode
R30842 N30841 N30842 10
D30842 N30842 0 diode
R30843 N30842 N30843 10
D30843 N30843 0 diode
R30844 N30843 N30844 10
D30844 N30844 0 diode
R30845 N30844 N30845 10
D30845 N30845 0 diode
R30846 N30845 N30846 10
D30846 N30846 0 diode
R30847 N30846 N30847 10
D30847 N30847 0 diode
R30848 N30847 N30848 10
D30848 N30848 0 diode
R30849 N30848 N30849 10
D30849 N30849 0 diode
R30850 N30849 N30850 10
D30850 N30850 0 diode
R30851 N30850 N30851 10
D30851 N30851 0 diode
R30852 N30851 N30852 10
D30852 N30852 0 diode
R30853 N30852 N30853 10
D30853 N30853 0 diode
R30854 N30853 N30854 10
D30854 N30854 0 diode
R30855 N30854 N30855 10
D30855 N30855 0 diode
R30856 N30855 N30856 10
D30856 N30856 0 diode
R30857 N30856 N30857 10
D30857 N30857 0 diode
R30858 N30857 N30858 10
D30858 N30858 0 diode
R30859 N30858 N30859 10
D30859 N30859 0 diode
R30860 N30859 N30860 10
D30860 N30860 0 diode
R30861 N30860 N30861 10
D30861 N30861 0 diode
R30862 N30861 N30862 10
D30862 N30862 0 diode
R30863 N30862 N30863 10
D30863 N30863 0 diode
R30864 N30863 N30864 10
D30864 N30864 0 diode
R30865 N30864 N30865 10
D30865 N30865 0 diode
R30866 N30865 N30866 10
D30866 N30866 0 diode
R30867 N30866 N30867 10
D30867 N30867 0 diode
R30868 N30867 N30868 10
D30868 N30868 0 diode
R30869 N30868 N30869 10
D30869 N30869 0 diode
R30870 N30869 N30870 10
D30870 N30870 0 diode
R30871 N30870 N30871 10
D30871 N30871 0 diode
R30872 N30871 N30872 10
D30872 N30872 0 diode
R30873 N30872 N30873 10
D30873 N30873 0 diode
R30874 N30873 N30874 10
D30874 N30874 0 diode
R30875 N30874 N30875 10
D30875 N30875 0 diode
R30876 N30875 N30876 10
D30876 N30876 0 diode
R30877 N30876 N30877 10
D30877 N30877 0 diode
R30878 N30877 N30878 10
D30878 N30878 0 diode
R30879 N30878 N30879 10
D30879 N30879 0 diode
R30880 N30879 N30880 10
D30880 N30880 0 diode
R30881 N30880 N30881 10
D30881 N30881 0 diode
R30882 N30881 N30882 10
D30882 N30882 0 diode
R30883 N30882 N30883 10
D30883 N30883 0 diode
R30884 N30883 N30884 10
D30884 N30884 0 diode
R30885 N30884 N30885 10
D30885 N30885 0 diode
R30886 N30885 N30886 10
D30886 N30886 0 diode
R30887 N30886 N30887 10
D30887 N30887 0 diode
R30888 N30887 N30888 10
D30888 N30888 0 diode
R30889 N30888 N30889 10
D30889 N30889 0 diode
R30890 N30889 N30890 10
D30890 N30890 0 diode
R30891 N30890 N30891 10
D30891 N30891 0 diode
R30892 N30891 N30892 10
D30892 N30892 0 diode
R30893 N30892 N30893 10
D30893 N30893 0 diode
R30894 N30893 N30894 10
D30894 N30894 0 diode
R30895 N30894 N30895 10
D30895 N30895 0 diode
R30896 N30895 N30896 10
D30896 N30896 0 diode
R30897 N30896 N30897 10
D30897 N30897 0 diode
R30898 N30897 N30898 10
D30898 N30898 0 diode
R30899 N30898 N30899 10
D30899 N30899 0 diode
R30900 N30899 N30900 10
D30900 N30900 0 diode
R30901 N30900 N30901 10
D30901 N30901 0 diode
R30902 N30901 N30902 10
D30902 N30902 0 diode
R30903 N30902 N30903 10
D30903 N30903 0 diode
R30904 N30903 N30904 10
D30904 N30904 0 diode
R30905 N30904 N30905 10
D30905 N30905 0 diode
R30906 N30905 N30906 10
D30906 N30906 0 diode
R30907 N30906 N30907 10
D30907 N30907 0 diode
R30908 N30907 N30908 10
D30908 N30908 0 diode
R30909 N30908 N30909 10
D30909 N30909 0 diode
R30910 N30909 N30910 10
D30910 N30910 0 diode
R30911 N30910 N30911 10
D30911 N30911 0 diode
R30912 N30911 N30912 10
D30912 N30912 0 diode
R30913 N30912 N30913 10
D30913 N30913 0 diode
R30914 N30913 N30914 10
D30914 N30914 0 diode
R30915 N30914 N30915 10
D30915 N30915 0 diode
R30916 N30915 N30916 10
D30916 N30916 0 diode
R30917 N30916 N30917 10
D30917 N30917 0 diode
R30918 N30917 N30918 10
D30918 N30918 0 diode
R30919 N30918 N30919 10
D30919 N30919 0 diode
R30920 N30919 N30920 10
D30920 N30920 0 diode
R30921 N30920 N30921 10
D30921 N30921 0 diode
R30922 N30921 N30922 10
D30922 N30922 0 diode
R30923 N30922 N30923 10
D30923 N30923 0 diode
R30924 N30923 N30924 10
D30924 N30924 0 diode
R30925 N30924 N30925 10
D30925 N30925 0 diode
R30926 N30925 N30926 10
D30926 N30926 0 diode
R30927 N30926 N30927 10
D30927 N30927 0 diode
R30928 N30927 N30928 10
D30928 N30928 0 diode
R30929 N30928 N30929 10
D30929 N30929 0 diode
R30930 N30929 N30930 10
D30930 N30930 0 diode
R30931 N30930 N30931 10
D30931 N30931 0 diode
R30932 N30931 N30932 10
D30932 N30932 0 diode
R30933 N30932 N30933 10
D30933 N30933 0 diode
R30934 N30933 N30934 10
D30934 N30934 0 diode
R30935 N30934 N30935 10
D30935 N30935 0 diode
R30936 N30935 N30936 10
D30936 N30936 0 diode
R30937 N30936 N30937 10
D30937 N30937 0 diode
R30938 N30937 N30938 10
D30938 N30938 0 diode
R30939 N30938 N30939 10
D30939 N30939 0 diode
R30940 N30939 N30940 10
D30940 N30940 0 diode
R30941 N30940 N30941 10
D30941 N30941 0 diode
R30942 N30941 N30942 10
D30942 N30942 0 diode
R30943 N30942 N30943 10
D30943 N30943 0 diode
R30944 N30943 N30944 10
D30944 N30944 0 diode
R30945 N30944 N30945 10
D30945 N30945 0 diode
R30946 N30945 N30946 10
D30946 N30946 0 diode
R30947 N30946 N30947 10
D30947 N30947 0 diode
R30948 N30947 N30948 10
D30948 N30948 0 diode
R30949 N30948 N30949 10
D30949 N30949 0 diode
R30950 N30949 N30950 10
D30950 N30950 0 diode
R30951 N30950 N30951 10
D30951 N30951 0 diode
R30952 N30951 N30952 10
D30952 N30952 0 diode
R30953 N30952 N30953 10
D30953 N30953 0 diode
R30954 N30953 N30954 10
D30954 N30954 0 diode
R30955 N30954 N30955 10
D30955 N30955 0 diode
R30956 N30955 N30956 10
D30956 N30956 0 diode
R30957 N30956 N30957 10
D30957 N30957 0 diode
R30958 N30957 N30958 10
D30958 N30958 0 diode
R30959 N30958 N30959 10
D30959 N30959 0 diode
R30960 N30959 N30960 10
D30960 N30960 0 diode
R30961 N30960 N30961 10
D30961 N30961 0 diode
R30962 N30961 N30962 10
D30962 N30962 0 diode
R30963 N30962 N30963 10
D30963 N30963 0 diode
R30964 N30963 N30964 10
D30964 N30964 0 diode
R30965 N30964 N30965 10
D30965 N30965 0 diode
R30966 N30965 N30966 10
D30966 N30966 0 diode
R30967 N30966 N30967 10
D30967 N30967 0 diode
R30968 N30967 N30968 10
D30968 N30968 0 diode
R30969 N30968 N30969 10
D30969 N30969 0 diode
R30970 N30969 N30970 10
D30970 N30970 0 diode
R30971 N30970 N30971 10
D30971 N30971 0 diode
R30972 N30971 N30972 10
D30972 N30972 0 diode
R30973 N30972 N30973 10
D30973 N30973 0 diode
R30974 N30973 N30974 10
D30974 N30974 0 diode
R30975 N30974 N30975 10
D30975 N30975 0 diode
R30976 N30975 N30976 10
D30976 N30976 0 diode
R30977 N30976 N30977 10
D30977 N30977 0 diode
R30978 N30977 N30978 10
D30978 N30978 0 diode
R30979 N30978 N30979 10
D30979 N30979 0 diode
R30980 N30979 N30980 10
D30980 N30980 0 diode
R30981 N30980 N30981 10
D30981 N30981 0 diode
R30982 N30981 N30982 10
D30982 N30982 0 diode
R30983 N30982 N30983 10
D30983 N30983 0 diode
R30984 N30983 N30984 10
D30984 N30984 0 diode
R30985 N30984 N30985 10
D30985 N30985 0 diode
R30986 N30985 N30986 10
D30986 N30986 0 diode
R30987 N30986 N30987 10
D30987 N30987 0 diode
R30988 N30987 N30988 10
D30988 N30988 0 diode
R30989 N30988 N30989 10
D30989 N30989 0 diode
R30990 N30989 N30990 10
D30990 N30990 0 diode
R30991 N30990 N30991 10
D30991 N30991 0 diode
R30992 N30991 N30992 10
D30992 N30992 0 diode
R30993 N30992 N30993 10
D30993 N30993 0 diode
R30994 N30993 N30994 10
D30994 N30994 0 diode
R30995 N30994 N30995 10
D30995 N30995 0 diode
R30996 N30995 N30996 10
D30996 N30996 0 diode
R30997 N30996 N30997 10
D30997 N30997 0 diode
R30998 N30997 N30998 10
D30998 N30998 0 diode
R30999 N30998 N30999 10
D30999 N30999 0 diode
R31000 N30999 N31000 10
D31000 N31000 0 diode
R31001 N31000 N31001 10
D31001 N31001 0 diode
R31002 N31001 N31002 10
D31002 N31002 0 diode
R31003 N31002 N31003 10
D31003 N31003 0 diode
R31004 N31003 N31004 10
D31004 N31004 0 diode
R31005 N31004 N31005 10
D31005 N31005 0 diode
R31006 N31005 N31006 10
D31006 N31006 0 diode
R31007 N31006 N31007 10
D31007 N31007 0 diode
R31008 N31007 N31008 10
D31008 N31008 0 diode
R31009 N31008 N31009 10
D31009 N31009 0 diode
R31010 N31009 N31010 10
D31010 N31010 0 diode
R31011 N31010 N31011 10
D31011 N31011 0 diode
R31012 N31011 N31012 10
D31012 N31012 0 diode
R31013 N31012 N31013 10
D31013 N31013 0 diode
R31014 N31013 N31014 10
D31014 N31014 0 diode
R31015 N31014 N31015 10
D31015 N31015 0 diode
R31016 N31015 N31016 10
D31016 N31016 0 diode
R31017 N31016 N31017 10
D31017 N31017 0 diode
R31018 N31017 N31018 10
D31018 N31018 0 diode
R31019 N31018 N31019 10
D31019 N31019 0 diode
R31020 N31019 N31020 10
D31020 N31020 0 diode
R31021 N31020 N31021 10
D31021 N31021 0 diode
R31022 N31021 N31022 10
D31022 N31022 0 diode
R31023 N31022 N31023 10
D31023 N31023 0 diode
R31024 N31023 N31024 10
D31024 N31024 0 diode
R31025 N31024 N31025 10
D31025 N31025 0 diode
R31026 N31025 N31026 10
D31026 N31026 0 diode
R31027 N31026 N31027 10
D31027 N31027 0 diode
R31028 N31027 N31028 10
D31028 N31028 0 diode
R31029 N31028 N31029 10
D31029 N31029 0 diode
R31030 N31029 N31030 10
D31030 N31030 0 diode
R31031 N31030 N31031 10
D31031 N31031 0 diode
R31032 N31031 N31032 10
D31032 N31032 0 diode
R31033 N31032 N31033 10
D31033 N31033 0 diode
R31034 N31033 N31034 10
D31034 N31034 0 diode
R31035 N31034 N31035 10
D31035 N31035 0 diode
R31036 N31035 N31036 10
D31036 N31036 0 diode
R31037 N31036 N31037 10
D31037 N31037 0 diode
R31038 N31037 N31038 10
D31038 N31038 0 diode
R31039 N31038 N31039 10
D31039 N31039 0 diode
R31040 N31039 N31040 10
D31040 N31040 0 diode
R31041 N31040 N31041 10
D31041 N31041 0 diode
R31042 N31041 N31042 10
D31042 N31042 0 diode
R31043 N31042 N31043 10
D31043 N31043 0 diode
R31044 N31043 N31044 10
D31044 N31044 0 diode
R31045 N31044 N31045 10
D31045 N31045 0 diode
R31046 N31045 N31046 10
D31046 N31046 0 diode
R31047 N31046 N31047 10
D31047 N31047 0 diode
R31048 N31047 N31048 10
D31048 N31048 0 diode
R31049 N31048 N31049 10
D31049 N31049 0 diode
R31050 N31049 N31050 10
D31050 N31050 0 diode
R31051 N31050 N31051 10
D31051 N31051 0 diode
R31052 N31051 N31052 10
D31052 N31052 0 diode
R31053 N31052 N31053 10
D31053 N31053 0 diode
R31054 N31053 N31054 10
D31054 N31054 0 diode
R31055 N31054 N31055 10
D31055 N31055 0 diode
R31056 N31055 N31056 10
D31056 N31056 0 diode
R31057 N31056 N31057 10
D31057 N31057 0 diode
R31058 N31057 N31058 10
D31058 N31058 0 diode
R31059 N31058 N31059 10
D31059 N31059 0 diode
R31060 N31059 N31060 10
D31060 N31060 0 diode
R31061 N31060 N31061 10
D31061 N31061 0 diode
R31062 N31061 N31062 10
D31062 N31062 0 diode
R31063 N31062 N31063 10
D31063 N31063 0 diode
R31064 N31063 N31064 10
D31064 N31064 0 diode
R31065 N31064 N31065 10
D31065 N31065 0 diode
R31066 N31065 N31066 10
D31066 N31066 0 diode
R31067 N31066 N31067 10
D31067 N31067 0 diode
R31068 N31067 N31068 10
D31068 N31068 0 diode
R31069 N31068 N31069 10
D31069 N31069 0 diode
R31070 N31069 N31070 10
D31070 N31070 0 diode
R31071 N31070 N31071 10
D31071 N31071 0 diode
R31072 N31071 N31072 10
D31072 N31072 0 diode
R31073 N31072 N31073 10
D31073 N31073 0 diode
R31074 N31073 N31074 10
D31074 N31074 0 diode
R31075 N31074 N31075 10
D31075 N31075 0 diode
R31076 N31075 N31076 10
D31076 N31076 0 diode
R31077 N31076 N31077 10
D31077 N31077 0 diode
R31078 N31077 N31078 10
D31078 N31078 0 diode
R31079 N31078 N31079 10
D31079 N31079 0 diode
R31080 N31079 N31080 10
D31080 N31080 0 diode
R31081 N31080 N31081 10
D31081 N31081 0 diode
R31082 N31081 N31082 10
D31082 N31082 0 diode
R31083 N31082 N31083 10
D31083 N31083 0 diode
R31084 N31083 N31084 10
D31084 N31084 0 diode
R31085 N31084 N31085 10
D31085 N31085 0 diode
R31086 N31085 N31086 10
D31086 N31086 0 diode
R31087 N31086 N31087 10
D31087 N31087 0 diode
R31088 N31087 N31088 10
D31088 N31088 0 diode
R31089 N31088 N31089 10
D31089 N31089 0 diode
R31090 N31089 N31090 10
D31090 N31090 0 diode
R31091 N31090 N31091 10
D31091 N31091 0 diode
R31092 N31091 N31092 10
D31092 N31092 0 diode
R31093 N31092 N31093 10
D31093 N31093 0 diode
R31094 N31093 N31094 10
D31094 N31094 0 diode
R31095 N31094 N31095 10
D31095 N31095 0 diode
R31096 N31095 N31096 10
D31096 N31096 0 diode
R31097 N31096 N31097 10
D31097 N31097 0 diode
R31098 N31097 N31098 10
D31098 N31098 0 diode
R31099 N31098 N31099 10
D31099 N31099 0 diode
R31100 N31099 N31100 10
D31100 N31100 0 diode
R31101 N31100 N31101 10
D31101 N31101 0 diode
R31102 N31101 N31102 10
D31102 N31102 0 diode
R31103 N31102 N31103 10
D31103 N31103 0 diode
R31104 N31103 N31104 10
D31104 N31104 0 diode
R31105 N31104 N31105 10
D31105 N31105 0 diode
R31106 N31105 N31106 10
D31106 N31106 0 diode
R31107 N31106 N31107 10
D31107 N31107 0 diode
R31108 N31107 N31108 10
D31108 N31108 0 diode
R31109 N31108 N31109 10
D31109 N31109 0 diode
R31110 N31109 N31110 10
D31110 N31110 0 diode
R31111 N31110 N31111 10
D31111 N31111 0 diode
R31112 N31111 N31112 10
D31112 N31112 0 diode
R31113 N31112 N31113 10
D31113 N31113 0 diode
R31114 N31113 N31114 10
D31114 N31114 0 diode
R31115 N31114 N31115 10
D31115 N31115 0 diode
R31116 N31115 N31116 10
D31116 N31116 0 diode
R31117 N31116 N31117 10
D31117 N31117 0 diode
R31118 N31117 N31118 10
D31118 N31118 0 diode
R31119 N31118 N31119 10
D31119 N31119 0 diode
R31120 N31119 N31120 10
D31120 N31120 0 diode
R31121 N31120 N31121 10
D31121 N31121 0 diode
R31122 N31121 N31122 10
D31122 N31122 0 diode
R31123 N31122 N31123 10
D31123 N31123 0 diode
R31124 N31123 N31124 10
D31124 N31124 0 diode
R31125 N31124 N31125 10
D31125 N31125 0 diode
R31126 N31125 N31126 10
D31126 N31126 0 diode
R31127 N31126 N31127 10
D31127 N31127 0 diode
R31128 N31127 N31128 10
D31128 N31128 0 diode
R31129 N31128 N31129 10
D31129 N31129 0 diode
R31130 N31129 N31130 10
D31130 N31130 0 diode
R31131 N31130 N31131 10
D31131 N31131 0 diode
R31132 N31131 N31132 10
D31132 N31132 0 diode
R31133 N31132 N31133 10
D31133 N31133 0 diode
R31134 N31133 N31134 10
D31134 N31134 0 diode
R31135 N31134 N31135 10
D31135 N31135 0 diode
R31136 N31135 N31136 10
D31136 N31136 0 diode
R31137 N31136 N31137 10
D31137 N31137 0 diode
R31138 N31137 N31138 10
D31138 N31138 0 diode
R31139 N31138 N31139 10
D31139 N31139 0 diode
R31140 N31139 N31140 10
D31140 N31140 0 diode
R31141 N31140 N31141 10
D31141 N31141 0 diode
R31142 N31141 N31142 10
D31142 N31142 0 diode
R31143 N31142 N31143 10
D31143 N31143 0 diode
R31144 N31143 N31144 10
D31144 N31144 0 diode
R31145 N31144 N31145 10
D31145 N31145 0 diode
R31146 N31145 N31146 10
D31146 N31146 0 diode
R31147 N31146 N31147 10
D31147 N31147 0 diode
R31148 N31147 N31148 10
D31148 N31148 0 diode
R31149 N31148 N31149 10
D31149 N31149 0 diode
R31150 N31149 N31150 10
D31150 N31150 0 diode
R31151 N31150 N31151 10
D31151 N31151 0 diode
R31152 N31151 N31152 10
D31152 N31152 0 diode
R31153 N31152 N31153 10
D31153 N31153 0 diode
R31154 N31153 N31154 10
D31154 N31154 0 diode
R31155 N31154 N31155 10
D31155 N31155 0 diode
R31156 N31155 N31156 10
D31156 N31156 0 diode
R31157 N31156 N31157 10
D31157 N31157 0 diode
R31158 N31157 N31158 10
D31158 N31158 0 diode
R31159 N31158 N31159 10
D31159 N31159 0 diode
R31160 N31159 N31160 10
D31160 N31160 0 diode
R31161 N31160 N31161 10
D31161 N31161 0 diode
R31162 N31161 N31162 10
D31162 N31162 0 diode
R31163 N31162 N31163 10
D31163 N31163 0 diode
R31164 N31163 N31164 10
D31164 N31164 0 diode
R31165 N31164 N31165 10
D31165 N31165 0 diode
R31166 N31165 N31166 10
D31166 N31166 0 diode
R31167 N31166 N31167 10
D31167 N31167 0 diode
R31168 N31167 N31168 10
D31168 N31168 0 diode
R31169 N31168 N31169 10
D31169 N31169 0 diode
R31170 N31169 N31170 10
D31170 N31170 0 diode
R31171 N31170 N31171 10
D31171 N31171 0 diode
R31172 N31171 N31172 10
D31172 N31172 0 diode
R31173 N31172 N31173 10
D31173 N31173 0 diode
R31174 N31173 N31174 10
D31174 N31174 0 diode
R31175 N31174 N31175 10
D31175 N31175 0 diode
R31176 N31175 N31176 10
D31176 N31176 0 diode
R31177 N31176 N31177 10
D31177 N31177 0 diode
R31178 N31177 N31178 10
D31178 N31178 0 diode
R31179 N31178 N31179 10
D31179 N31179 0 diode
R31180 N31179 N31180 10
D31180 N31180 0 diode
R31181 N31180 N31181 10
D31181 N31181 0 diode
R31182 N31181 N31182 10
D31182 N31182 0 diode
R31183 N31182 N31183 10
D31183 N31183 0 diode
R31184 N31183 N31184 10
D31184 N31184 0 diode
R31185 N31184 N31185 10
D31185 N31185 0 diode
R31186 N31185 N31186 10
D31186 N31186 0 diode
R31187 N31186 N31187 10
D31187 N31187 0 diode
R31188 N31187 N31188 10
D31188 N31188 0 diode
R31189 N31188 N31189 10
D31189 N31189 0 diode
R31190 N31189 N31190 10
D31190 N31190 0 diode
R31191 N31190 N31191 10
D31191 N31191 0 diode
R31192 N31191 N31192 10
D31192 N31192 0 diode
R31193 N31192 N31193 10
D31193 N31193 0 diode
R31194 N31193 N31194 10
D31194 N31194 0 diode
R31195 N31194 N31195 10
D31195 N31195 0 diode
R31196 N31195 N31196 10
D31196 N31196 0 diode
R31197 N31196 N31197 10
D31197 N31197 0 diode
R31198 N31197 N31198 10
D31198 N31198 0 diode
R31199 N31198 N31199 10
D31199 N31199 0 diode
R31200 N31199 N31200 10
D31200 N31200 0 diode
R31201 N31200 N31201 10
D31201 N31201 0 diode
R31202 N31201 N31202 10
D31202 N31202 0 diode
R31203 N31202 N31203 10
D31203 N31203 0 diode
R31204 N31203 N31204 10
D31204 N31204 0 diode
R31205 N31204 N31205 10
D31205 N31205 0 diode
R31206 N31205 N31206 10
D31206 N31206 0 diode
R31207 N31206 N31207 10
D31207 N31207 0 diode
R31208 N31207 N31208 10
D31208 N31208 0 diode
R31209 N31208 N31209 10
D31209 N31209 0 diode
R31210 N31209 N31210 10
D31210 N31210 0 diode
R31211 N31210 N31211 10
D31211 N31211 0 diode
R31212 N31211 N31212 10
D31212 N31212 0 diode
R31213 N31212 N31213 10
D31213 N31213 0 diode
R31214 N31213 N31214 10
D31214 N31214 0 diode
R31215 N31214 N31215 10
D31215 N31215 0 diode
R31216 N31215 N31216 10
D31216 N31216 0 diode
R31217 N31216 N31217 10
D31217 N31217 0 diode
R31218 N31217 N31218 10
D31218 N31218 0 diode
R31219 N31218 N31219 10
D31219 N31219 0 diode
R31220 N31219 N31220 10
D31220 N31220 0 diode
R31221 N31220 N31221 10
D31221 N31221 0 diode
R31222 N31221 N31222 10
D31222 N31222 0 diode
R31223 N31222 N31223 10
D31223 N31223 0 diode
R31224 N31223 N31224 10
D31224 N31224 0 diode
R31225 N31224 N31225 10
D31225 N31225 0 diode
R31226 N31225 N31226 10
D31226 N31226 0 diode
R31227 N31226 N31227 10
D31227 N31227 0 diode
R31228 N31227 N31228 10
D31228 N31228 0 diode
R31229 N31228 N31229 10
D31229 N31229 0 diode
R31230 N31229 N31230 10
D31230 N31230 0 diode
R31231 N31230 N31231 10
D31231 N31231 0 diode
R31232 N31231 N31232 10
D31232 N31232 0 diode
R31233 N31232 N31233 10
D31233 N31233 0 diode
R31234 N31233 N31234 10
D31234 N31234 0 diode
R31235 N31234 N31235 10
D31235 N31235 0 diode
R31236 N31235 N31236 10
D31236 N31236 0 diode
R31237 N31236 N31237 10
D31237 N31237 0 diode
R31238 N31237 N31238 10
D31238 N31238 0 diode
R31239 N31238 N31239 10
D31239 N31239 0 diode
R31240 N31239 N31240 10
D31240 N31240 0 diode
R31241 N31240 N31241 10
D31241 N31241 0 diode
R31242 N31241 N31242 10
D31242 N31242 0 diode
R31243 N31242 N31243 10
D31243 N31243 0 diode
R31244 N31243 N31244 10
D31244 N31244 0 diode
R31245 N31244 N31245 10
D31245 N31245 0 diode
R31246 N31245 N31246 10
D31246 N31246 0 diode
R31247 N31246 N31247 10
D31247 N31247 0 diode
R31248 N31247 N31248 10
D31248 N31248 0 diode
R31249 N31248 N31249 10
D31249 N31249 0 diode
R31250 N31249 N31250 10
D31250 N31250 0 diode
R31251 N31250 N31251 10
D31251 N31251 0 diode
R31252 N31251 N31252 10
D31252 N31252 0 diode
R31253 N31252 N31253 10
D31253 N31253 0 diode
R31254 N31253 N31254 10
D31254 N31254 0 diode
R31255 N31254 N31255 10
D31255 N31255 0 diode
R31256 N31255 N31256 10
D31256 N31256 0 diode
R31257 N31256 N31257 10
D31257 N31257 0 diode
R31258 N31257 N31258 10
D31258 N31258 0 diode
R31259 N31258 N31259 10
D31259 N31259 0 diode
R31260 N31259 N31260 10
D31260 N31260 0 diode
R31261 N31260 N31261 10
D31261 N31261 0 diode
R31262 N31261 N31262 10
D31262 N31262 0 diode
R31263 N31262 N31263 10
D31263 N31263 0 diode
R31264 N31263 N31264 10
D31264 N31264 0 diode
R31265 N31264 N31265 10
D31265 N31265 0 diode
R31266 N31265 N31266 10
D31266 N31266 0 diode
R31267 N31266 N31267 10
D31267 N31267 0 diode
R31268 N31267 N31268 10
D31268 N31268 0 diode
R31269 N31268 N31269 10
D31269 N31269 0 diode
R31270 N31269 N31270 10
D31270 N31270 0 diode
R31271 N31270 N31271 10
D31271 N31271 0 diode
R31272 N31271 N31272 10
D31272 N31272 0 diode
R31273 N31272 N31273 10
D31273 N31273 0 diode
R31274 N31273 N31274 10
D31274 N31274 0 diode
R31275 N31274 N31275 10
D31275 N31275 0 diode
R31276 N31275 N31276 10
D31276 N31276 0 diode
R31277 N31276 N31277 10
D31277 N31277 0 diode
R31278 N31277 N31278 10
D31278 N31278 0 diode
R31279 N31278 N31279 10
D31279 N31279 0 diode
R31280 N31279 N31280 10
D31280 N31280 0 diode
R31281 N31280 N31281 10
D31281 N31281 0 diode
R31282 N31281 N31282 10
D31282 N31282 0 diode
R31283 N31282 N31283 10
D31283 N31283 0 diode
R31284 N31283 N31284 10
D31284 N31284 0 diode
R31285 N31284 N31285 10
D31285 N31285 0 diode
R31286 N31285 N31286 10
D31286 N31286 0 diode
R31287 N31286 N31287 10
D31287 N31287 0 diode
R31288 N31287 N31288 10
D31288 N31288 0 diode
R31289 N31288 N31289 10
D31289 N31289 0 diode
R31290 N31289 N31290 10
D31290 N31290 0 diode
R31291 N31290 N31291 10
D31291 N31291 0 diode
R31292 N31291 N31292 10
D31292 N31292 0 diode
R31293 N31292 N31293 10
D31293 N31293 0 diode
R31294 N31293 N31294 10
D31294 N31294 0 diode
R31295 N31294 N31295 10
D31295 N31295 0 diode
R31296 N31295 N31296 10
D31296 N31296 0 diode
R31297 N31296 N31297 10
D31297 N31297 0 diode
R31298 N31297 N31298 10
D31298 N31298 0 diode
R31299 N31298 N31299 10
D31299 N31299 0 diode
R31300 N31299 N31300 10
D31300 N31300 0 diode
R31301 N31300 N31301 10
D31301 N31301 0 diode
R31302 N31301 N31302 10
D31302 N31302 0 diode
R31303 N31302 N31303 10
D31303 N31303 0 diode
R31304 N31303 N31304 10
D31304 N31304 0 diode
R31305 N31304 N31305 10
D31305 N31305 0 diode
R31306 N31305 N31306 10
D31306 N31306 0 diode
R31307 N31306 N31307 10
D31307 N31307 0 diode
R31308 N31307 N31308 10
D31308 N31308 0 diode
R31309 N31308 N31309 10
D31309 N31309 0 diode
R31310 N31309 N31310 10
D31310 N31310 0 diode
R31311 N31310 N31311 10
D31311 N31311 0 diode
R31312 N31311 N31312 10
D31312 N31312 0 diode
R31313 N31312 N31313 10
D31313 N31313 0 diode
R31314 N31313 N31314 10
D31314 N31314 0 diode
R31315 N31314 N31315 10
D31315 N31315 0 diode
R31316 N31315 N31316 10
D31316 N31316 0 diode
R31317 N31316 N31317 10
D31317 N31317 0 diode
R31318 N31317 N31318 10
D31318 N31318 0 diode
R31319 N31318 N31319 10
D31319 N31319 0 diode
R31320 N31319 N31320 10
D31320 N31320 0 diode
R31321 N31320 N31321 10
D31321 N31321 0 diode
R31322 N31321 N31322 10
D31322 N31322 0 diode
R31323 N31322 N31323 10
D31323 N31323 0 diode
R31324 N31323 N31324 10
D31324 N31324 0 diode
R31325 N31324 N31325 10
D31325 N31325 0 diode
R31326 N31325 N31326 10
D31326 N31326 0 diode
R31327 N31326 N31327 10
D31327 N31327 0 diode
R31328 N31327 N31328 10
D31328 N31328 0 diode
R31329 N31328 N31329 10
D31329 N31329 0 diode
R31330 N31329 N31330 10
D31330 N31330 0 diode
R31331 N31330 N31331 10
D31331 N31331 0 diode
R31332 N31331 N31332 10
D31332 N31332 0 diode
R31333 N31332 N31333 10
D31333 N31333 0 diode
R31334 N31333 N31334 10
D31334 N31334 0 diode
R31335 N31334 N31335 10
D31335 N31335 0 diode
R31336 N31335 N31336 10
D31336 N31336 0 diode
R31337 N31336 N31337 10
D31337 N31337 0 diode
R31338 N31337 N31338 10
D31338 N31338 0 diode
R31339 N31338 N31339 10
D31339 N31339 0 diode
R31340 N31339 N31340 10
D31340 N31340 0 diode
R31341 N31340 N31341 10
D31341 N31341 0 diode
R31342 N31341 N31342 10
D31342 N31342 0 diode
R31343 N31342 N31343 10
D31343 N31343 0 diode
R31344 N31343 N31344 10
D31344 N31344 0 diode
R31345 N31344 N31345 10
D31345 N31345 0 diode
R31346 N31345 N31346 10
D31346 N31346 0 diode
R31347 N31346 N31347 10
D31347 N31347 0 diode
R31348 N31347 N31348 10
D31348 N31348 0 diode
R31349 N31348 N31349 10
D31349 N31349 0 diode
R31350 N31349 N31350 10
D31350 N31350 0 diode
R31351 N31350 N31351 10
D31351 N31351 0 diode
R31352 N31351 N31352 10
D31352 N31352 0 diode
R31353 N31352 N31353 10
D31353 N31353 0 diode
R31354 N31353 N31354 10
D31354 N31354 0 diode
R31355 N31354 N31355 10
D31355 N31355 0 diode
R31356 N31355 N31356 10
D31356 N31356 0 diode
R31357 N31356 N31357 10
D31357 N31357 0 diode
R31358 N31357 N31358 10
D31358 N31358 0 diode
R31359 N31358 N31359 10
D31359 N31359 0 diode
R31360 N31359 N31360 10
D31360 N31360 0 diode
R31361 N31360 N31361 10
D31361 N31361 0 diode
R31362 N31361 N31362 10
D31362 N31362 0 diode
R31363 N31362 N31363 10
D31363 N31363 0 diode
R31364 N31363 N31364 10
D31364 N31364 0 diode
R31365 N31364 N31365 10
D31365 N31365 0 diode
R31366 N31365 N31366 10
D31366 N31366 0 diode
R31367 N31366 N31367 10
D31367 N31367 0 diode
R31368 N31367 N31368 10
D31368 N31368 0 diode
R31369 N31368 N31369 10
D31369 N31369 0 diode
R31370 N31369 N31370 10
D31370 N31370 0 diode
R31371 N31370 N31371 10
D31371 N31371 0 diode
R31372 N31371 N31372 10
D31372 N31372 0 diode
R31373 N31372 N31373 10
D31373 N31373 0 diode
R31374 N31373 N31374 10
D31374 N31374 0 diode
R31375 N31374 N31375 10
D31375 N31375 0 diode
R31376 N31375 N31376 10
D31376 N31376 0 diode
R31377 N31376 N31377 10
D31377 N31377 0 diode
R31378 N31377 N31378 10
D31378 N31378 0 diode
R31379 N31378 N31379 10
D31379 N31379 0 diode
R31380 N31379 N31380 10
D31380 N31380 0 diode
R31381 N31380 N31381 10
D31381 N31381 0 diode
R31382 N31381 N31382 10
D31382 N31382 0 diode
R31383 N31382 N31383 10
D31383 N31383 0 diode
R31384 N31383 N31384 10
D31384 N31384 0 diode
R31385 N31384 N31385 10
D31385 N31385 0 diode
R31386 N31385 N31386 10
D31386 N31386 0 diode
R31387 N31386 N31387 10
D31387 N31387 0 diode
R31388 N31387 N31388 10
D31388 N31388 0 diode
R31389 N31388 N31389 10
D31389 N31389 0 diode
R31390 N31389 N31390 10
D31390 N31390 0 diode
R31391 N31390 N31391 10
D31391 N31391 0 diode
R31392 N31391 N31392 10
D31392 N31392 0 diode
R31393 N31392 N31393 10
D31393 N31393 0 diode
R31394 N31393 N31394 10
D31394 N31394 0 diode
R31395 N31394 N31395 10
D31395 N31395 0 diode
R31396 N31395 N31396 10
D31396 N31396 0 diode
R31397 N31396 N31397 10
D31397 N31397 0 diode
R31398 N31397 N31398 10
D31398 N31398 0 diode
R31399 N31398 N31399 10
D31399 N31399 0 diode
R31400 N31399 N31400 10
D31400 N31400 0 diode
R31401 N31400 N31401 10
D31401 N31401 0 diode
R31402 N31401 N31402 10
D31402 N31402 0 diode
R31403 N31402 N31403 10
D31403 N31403 0 diode
R31404 N31403 N31404 10
D31404 N31404 0 diode
R31405 N31404 N31405 10
D31405 N31405 0 diode
R31406 N31405 N31406 10
D31406 N31406 0 diode
R31407 N31406 N31407 10
D31407 N31407 0 diode
R31408 N31407 N31408 10
D31408 N31408 0 diode
R31409 N31408 N31409 10
D31409 N31409 0 diode
R31410 N31409 N31410 10
D31410 N31410 0 diode
R31411 N31410 N31411 10
D31411 N31411 0 diode
R31412 N31411 N31412 10
D31412 N31412 0 diode
R31413 N31412 N31413 10
D31413 N31413 0 diode
R31414 N31413 N31414 10
D31414 N31414 0 diode
R31415 N31414 N31415 10
D31415 N31415 0 diode
R31416 N31415 N31416 10
D31416 N31416 0 diode
R31417 N31416 N31417 10
D31417 N31417 0 diode
R31418 N31417 N31418 10
D31418 N31418 0 diode
R31419 N31418 N31419 10
D31419 N31419 0 diode
R31420 N31419 N31420 10
D31420 N31420 0 diode
R31421 N31420 N31421 10
D31421 N31421 0 diode
R31422 N31421 N31422 10
D31422 N31422 0 diode
R31423 N31422 N31423 10
D31423 N31423 0 diode
R31424 N31423 N31424 10
D31424 N31424 0 diode
R31425 N31424 N31425 10
D31425 N31425 0 diode
R31426 N31425 N31426 10
D31426 N31426 0 diode
R31427 N31426 N31427 10
D31427 N31427 0 diode
R31428 N31427 N31428 10
D31428 N31428 0 diode
R31429 N31428 N31429 10
D31429 N31429 0 diode
R31430 N31429 N31430 10
D31430 N31430 0 diode
R31431 N31430 N31431 10
D31431 N31431 0 diode
R31432 N31431 N31432 10
D31432 N31432 0 diode
R31433 N31432 N31433 10
D31433 N31433 0 diode
R31434 N31433 N31434 10
D31434 N31434 0 diode
R31435 N31434 N31435 10
D31435 N31435 0 diode
R31436 N31435 N31436 10
D31436 N31436 0 diode
R31437 N31436 N31437 10
D31437 N31437 0 diode
R31438 N31437 N31438 10
D31438 N31438 0 diode
R31439 N31438 N31439 10
D31439 N31439 0 diode
R31440 N31439 N31440 10
D31440 N31440 0 diode
R31441 N31440 N31441 10
D31441 N31441 0 diode
R31442 N31441 N31442 10
D31442 N31442 0 diode
R31443 N31442 N31443 10
D31443 N31443 0 diode
R31444 N31443 N31444 10
D31444 N31444 0 diode
R31445 N31444 N31445 10
D31445 N31445 0 diode
R31446 N31445 N31446 10
D31446 N31446 0 diode
R31447 N31446 N31447 10
D31447 N31447 0 diode
R31448 N31447 N31448 10
D31448 N31448 0 diode
R31449 N31448 N31449 10
D31449 N31449 0 diode
R31450 N31449 N31450 10
D31450 N31450 0 diode
R31451 N31450 N31451 10
D31451 N31451 0 diode
R31452 N31451 N31452 10
D31452 N31452 0 diode
R31453 N31452 N31453 10
D31453 N31453 0 diode
R31454 N31453 N31454 10
D31454 N31454 0 diode
R31455 N31454 N31455 10
D31455 N31455 0 diode
R31456 N31455 N31456 10
D31456 N31456 0 diode
R31457 N31456 N31457 10
D31457 N31457 0 diode
R31458 N31457 N31458 10
D31458 N31458 0 diode
R31459 N31458 N31459 10
D31459 N31459 0 diode
R31460 N31459 N31460 10
D31460 N31460 0 diode
R31461 N31460 N31461 10
D31461 N31461 0 diode
R31462 N31461 N31462 10
D31462 N31462 0 diode
R31463 N31462 N31463 10
D31463 N31463 0 diode
R31464 N31463 N31464 10
D31464 N31464 0 diode
R31465 N31464 N31465 10
D31465 N31465 0 diode
R31466 N31465 N31466 10
D31466 N31466 0 diode
R31467 N31466 N31467 10
D31467 N31467 0 diode
R31468 N31467 N31468 10
D31468 N31468 0 diode
R31469 N31468 N31469 10
D31469 N31469 0 diode
R31470 N31469 N31470 10
D31470 N31470 0 diode
R31471 N31470 N31471 10
D31471 N31471 0 diode
R31472 N31471 N31472 10
D31472 N31472 0 diode
R31473 N31472 N31473 10
D31473 N31473 0 diode
R31474 N31473 N31474 10
D31474 N31474 0 diode
R31475 N31474 N31475 10
D31475 N31475 0 diode
R31476 N31475 N31476 10
D31476 N31476 0 diode
R31477 N31476 N31477 10
D31477 N31477 0 diode
R31478 N31477 N31478 10
D31478 N31478 0 diode
R31479 N31478 N31479 10
D31479 N31479 0 diode
R31480 N31479 N31480 10
D31480 N31480 0 diode
R31481 N31480 N31481 10
D31481 N31481 0 diode
R31482 N31481 N31482 10
D31482 N31482 0 diode
R31483 N31482 N31483 10
D31483 N31483 0 diode
R31484 N31483 N31484 10
D31484 N31484 0 diode
R31485 N31484 N31485 10
D31485 N31485 0 diode
R31486 N31485 N31486 10
D31486 N31486 0 diode
R31487 N31486 N31487 10
D31487 N31487 0 diode
R31488 N31487 N31488 10
D31488 N31488 0 diode
R31489 N31488 N31489 10
D31489 N31489 0 diode
R31490 N31489 N31490 10
D31490 N31490 0 diode
R31491 N31490 N31491 10
D31491 N31491 0 diode
R31492 N31491 N31492 10
D31492 N31492 0 diode
R31493 N31492 N31493 10
D31493 N31493 0 diode
R31494 N31493 N31494 10
D31494 N31494 0 diode
R31495 N31494 N31495 10
D31495 N31495 0 diode
R31496 N31495 N31496 10
D31496 N31496 0 diode
R31497 N31496 N31497 10
D31497 N31497 0 diode
R31498 N31497 N31498 10
D31498 N31498 0 diode
R31499 N31498 N31499 10
D31499 N31499 0 diode
R31500 N31499 N31500 10
D31500 N31500 0 diode
R31501 N31500 N31501 10
D31501 N31501 0 diode
R31502 N31501 N31502 10
D31502 N31502 0 diode
R31503 N31502 N31503 10
D31503 N31503 0 diode
R31504 N31503 N31504 10
D31504 N31504 0 diode
R31505 N31504 N31505 10
D31505 N31505 0 diode
R31506 N31505 N31506 10
D31506 N31506 0 diode
R31507 N31506 N31507 10
D31507 N31507 0 diode
R31508 N31507 N31508 10
D31508 N31508 0 diode
R31509 N31508 N31509 10
D31509 N31509 0 diode
R31510 N31509 N31510 10
D31510 N31510 0 diode
R31511 N31510 N31511 10
D31511 N31511 0 diode
R31512 N31511 N31512 10
D31512 N31512 0 diode
R31513 N31512 N31513 10
D31513 N31513 0 diode
R31514 N31513 N31514 10
D31514 N31514 0 diode
R31515 N31514 N31515 10
D31515 N31515 0 diode
R31516 N31515 N31516 10
D31516 N31516 0 diode
R31517 N31516 N31517 10
D31517 N31517 0 diode
R31518 N31517 N31518 10
D31518 N31518 0 diode
R31519 N31518 N31519 10
D31519 N31519 0 diode
R31520 N31519 N31520 10
D31520 N31520 0 diode
R31521 N31520 N31521 10
D31521 N31521 0 diode
R31522 N31521 N31522 10
D31522 N31522 0 diode
R31523 N31522 N31523 10
D31523 N31523 0 diode
R31524 N31523 N31524 10
D31524 N31524 0 diode
R31525 N31524 N31525 10
D31525 N31525 0 diode
R31526 N31525 N31526 10
D31526 N31526 0 diode
R31527 N31526 N31527 10
D31527 N31527 0 diode
R31528 N31527 N31528 10
D31528 N31528 0 diode
R31529 N31528 N31529 10
D31529 N31529 0 diode
R31530 N31529 N31530 10
D31530 N31530 0 diode
R31531 N31530 N31531 10
D31531 N31531 0 diode
R31532 N31531 N31532 10
D31532 N31532 0 diode
R31533 N31532 N31533 10
D31533 N31533 0 diode
R31534 N31533 N31534 10
D31534 N31534 0 diode
R31535 N31534 N31535 10
D31535 N31535 0 diode
R31536 N31535 N31536 10
D31536 N31536 0 diode
R31537 N31536 N31537 10
D31537 N31537 0 diode
R31538 N31537 N31538 10
D31538 N31538 0 diode
R31539 N31538 N31539 10
D31539 N31539 0 diode
R31540 N31539 N31540 10
D31540 N31540 0 diode
R31541 N31540 N31541 10
D31541 N31541 0 diode
R31542 N31541 N31542 10
D31542 N31542 0 diode
R31543 N31542 N31543 10
D31543 N31543 0 diode
R31544 N31543 N31544 10
D31544 N31544 0 diode
R31545 N31544 N31545 10
D31545 N31545 0 diode
R31546 N31545 N31546 10
D31546 N31546 0 diode
R31547 N31546 N31547 10
D31547 N31547 0 diode
R31548 N31547 N31548 10
D31548 N31548 0 diode
R31549 N31548 N31549 10
D31549 N31549 0 diode
R31550 N31549 N31550 10
D31550 N31550 0 diode
R31551 N31550 N31551 10
D31551 N31551 0 diode
R31552 N31551 N31552 10
D31552 N31552 0 diode
R31553 N31552 N31553 10
D31553 N31553 0 diode
R31554 N31553 N31554 10
D31554 N31554 0 diode
R31555 N31554 N31555 10
D31555 N31555 0 diode
R31556 N31555 N31556 10
D31556 N31556 0 diode
R31557 N31556 N31557 10
D31557 N31557 0 diode
R31558 N31557 N31558 10
D31558 N31558 0 diode
R31559 N31558 N31559 10
D31559 N31559 0 diode
R31560 N31559 N31560 10
D31560 N31560 0 diode
R31561 N31560 N31561 10
D31561 N31561 0 diode
R31562 N31561 N31562 10
D31562 N31562 0 diode
R31563 N31562 N31563 10
D31563 N31563 0 diode
R31564 N31563 N31564 10
D31564 N31564 0 diode
R31565 N31564 N31565 10
D31565 N31565 0 diode
R31566 N31565 N31566 10
D31566 N31566 0 diode
R31567 N31566 N31567 10
D31567 N31567 0 diode
R31568 N31567 N31568 10
D31568 N31568 0 diode
R31569 N31568 N31569 10
D31569 N31569 0 diode
R31570 N31569 N31570 10
D31570 N31570 0 diode
R31571 N31570 N31571 10
D31571 N31571 0 diode
R31572 N31571 N31572 10
D31572 N31572 0 diode
R31573 N31572 N31573 10
D31573 N31573 0 diode
R31574 N31573 N31574 10
D31574 N31574 0 diode
R31575 N31574 N31575 10
D31575 N31575 0 diode
R31576 N31575 N31576 10
D31576 N31576 0 diode
R31577 N31576 N31577 10
D31577 N31577 0 diode
R31578 N31577 N31578 10
D31578 N31578 0 diode
R31579 N31578 N31579 10
D31579 N31579 0 diode
R31580 N31579 N31580 10
D31580 N31580 0 diode
R31581 N31580 N31581 10
D31581 N31581 0 diode
R31582 N31581 N31582 10
D31582 N31582 0 diode
R31583 N31582 N31583 10
D31583 N31583 0 diode
R31584 N31583 N31584 10
D31584 N31584 0 diode
R31585 N31584 N31585 10
D31585 N31585 0 diode
R31586 N31585 N31586 10
D31586 N31586 0 diode
R31587 N31586 N31587 10
D31587 N31587 0 diode
R31588 N31587 N31588 10
D31588 N31588 0 diode
R31589 N31588 N31589 10
D31589 N31589 0 diode
R31590 N31589 N31590 10
D31590 N31590 0 diode
R31591 N31590 N31591 10
D31591 N31591 0 diode
R31592 N31591 N31592 10
D31592 N31592 0 diode
R31593 N31592 N31593 10
D31593 N31593 0 diode
R31594 N31593 N31594 10
D31594 N31594 0 diode
R31595 N31594 N31595 10
D31595 N31595 0 diode
R31596 N31595 N31596 10
D31596 N31596 0 diode
R31597 N31596 N31597 10
D31597 N31597 0 diode
R31598 N31597 N31598 10
D31598 N31598 0 diode
R31599 N31598 N31599 10
D31599 N31599 0 diode
R31600 N31599 N31600 10
D31600 N31600 0 diode
R31601 N31600 N31601 10
D31601 N31601 0 diode
R31602 N31601 N31602 10
D31602 N31602 0 diode
R31603 N31602 N31603 10
D31603 N31603 0 diode
R31604 N31603 N31604 10
D31604 N31604 0 diode
R31605 N31604 N31605 10
D31605 N31605 0 diode
R31606 N31605 N31606 10
D31606 N31606 0 diode
R31607 N31606 N31607 10
D31607 N31607 0 diode
R31608 N31607 N31608 10
D31608 N31608 0 diode
R31609 N31608 N31609 10
D31609 N31609 0 diode
R31610 N31609 N31610 10
D31610 N31610 0 diode
R31611 N31610 N31611 10
D31611 N31611 0 diode
R31612 N31611 N31612 10
D31612 N31612 0 diode
R31613 N31612 N31613 10
D31613 N31613 0 diode
R31614 N31613 N31614 10
D31614 N31614 0 diode
R31615 N31614 N31615 10
D31615 N31615 0 diode
R31616 N31615 N31616 10
D31616 N31616 0 diode
R31617 N31616 N31617 10
D31617 N31617 0 diode
R31618 N31617 N31618 10
D31618 N31618 0 diode
R31619 N31618 N31619 10
D31619 N31619 0 diode
R31620 N31619 N31620 10
D31620 N31620 0 diode
R31621 N31620 N31621 10
D31621 N31621 0 diode
R31622 N31621 N31622 10
D31622 N31622 0 diode
R31623 N31622 N31623 10
D31623 N31623 0 diode
R31624 N31623 N31624 10
D31624 N31624 0 diode
R31625 N31624 N31625 10
D31625 N31625 0 diode
R31626 N31625 N31626 10
D31626 N31626 0 diode
R31627 N31626 N31627 10
D31627 N31627 0 diode
R31628 N31627 N31628 10
D31628 N31628 0 diode
R31629 N31628 N31629 10
D31629 N31629 0 diode
R31630 N31629 N31630 10
D31630 N31630 0 diode
R31631 N31630 N31631 10
D31631 N31631 0 diode
R31632 N31631 N31632 10
D31632 N31632 0 diode
R31633 N31632 N31633 10
D31633 N31633 0 diode
R31634 N31633 N31634 10
D31634 N31634 0 diode
R31635 N31634 N31635 10
D31635 N31635 0 diode
R31636 N31635 N31636 10
D31636 N31636 0 diode
R31637 N31636 N31637 10
D31637 N31637 0 diode
R31638 N31637 N31638 10
D31638 N31638 0 diode
R31639 N31638 N31639 10
D31639 N31639 0 diode
R31640 N31639 N31640 10
D31640 N31640 0 diode
R31641 N31640 N31641 10
D31641 N31641 0 diode
R31642 N31641 N31642 10
D31642 N31642 0 diode
R31643 N31642 N31643 10
D31643 N31643 0 diode
R31644 N31643 N31644 10
D31644 N31644 0 diode
R31645 N31644 N31645 10
D31645 N31645 0 diode
R31646 N31645 N31646 10
D31646 N31646 0 diode
R31647 N31646 N31647 10
D31647 N31647 0 diode
R31648 N31647 N31648 10
D31648 N31648 0 diode
R31649 N31648 N31649 10
D31649 N31649 0 diode
R31650 N31649 N31650 10
D31650 N31650 0 diode
R31651 N31650 N31651 10
D31651 N31651 0 diode
R31652 N31651 N31652 10
D31652 N31652 0 diode
R31653 N31652 N31653 10
D31653 N31653 0 diode
R31654 N31653 N31654 10
D31654 N31654 0 diode
R31655 N31654 N31655 10
D31655 N31655 0 diode
R31656 N31655 N31656 10
D31656 N31656 0 diode
R31657 N31656 N31657 10
D31657 N31657 0 diode
R31658 N31657 N31658 10
D31658 N31658 0 diode
R31659 N31658 N31659 10
D31659 N31659 0 diode
R31660 N31659 N31660 10
D31660 N31660 0 diode
R31661 N31660 N31661 10
D31661 N31661 0 diode
R31662 N31661 N31662 10
D31662 N31662 0 diode
R31663 N31662 N31663 10
D31663 N31663 0 diode
R31664 N31663 N31664 10
D31664 N31664 0 diode
R31665 N31664 N31665 10
D31665 N31665 0 diode
R31666 N31665 N31666 10
D31666 N31666 0 diode
R31667 N31666 N31667 10
D31667 N31667 0 diode
R31668 N31667 N31668 10
D31668 N31668 0 diode
R31669 N31668 N31669 10
D31669 N31669 0 diode
R31670 N31669 N31670 10
D31670 N31670 0 diode
R31671 N31670 N31671 10
D31671 N31671 0 diode
R31672 N31671 N31672 10
D31672 N31672 0 diode
R31673 N31672 N31673 10
D31673 N31673 0 diode
R31674 N31673 N31674 10
D31674 N31674 0 diode
R31675 N31674 N31675 10
D31675 N31675 0 diode
R31676 N31675 N31676 10
D31676 N31676 0 diode
R31677 N31676 N31677 10
D31677 N31677 0 diode
R31678 N31677 N31678 10
D31678 N31678 0 diode
R31679 N31678 N31679 10
D31679 N31679 0 diode
R31680 N31679 N31680 10
D31680 N31680 0 diode
R31681 N31680 N31681 10
D31681 N31681 0 diode
R31682 N31681 N31682 10
D31682 N31682 0 diode
R31683 N31682 N31683 10
D31683 N31683 0 diode
R31684 N31683 N31684 10
D31684 N31684 0 diode
R31685 N31684 N31685 10
D31685 N31685 0 diode
R31686 N31685 N31686 10
D31686 N31686 0 diode
R31687 N31686 N31687 10
D31687 N31687 0 diode
R31688 N31687 N31688 10
D31688 N31688 0 diode
R31689 N31688 N31689 10
D31689 N31689 0 diode
R31690 N31689 N31690 10
D31690 N31690 0 diode
R31691 N31690 N31691 10
D31691 N31691 0 diode
R31692 N31691 N31692 10
D31692 N31692 0 diode
R31693 N31692 N31693 10
D31693 N31693 0 diode
R31694 N31693 N31694 10
D31694 N31694 0 diode
R31695 N31694 N31695 10
D31695 N31695 0 diode
R31696 N31695 N31696 10
D31696 N31696 0 diode
R31697 N31696 N31697 10
D31697 N31697 0 diode
R31698 N31697 N31698 10
D31698 N31698 0 diode
R31699 N31698 N31699 10
D31699 N31699 0 diode
R31700 N31699 N31700 10
D31700 N31700 0 diode
R31701 N31700 N31701 10
D31701 N31701 0 diode
R31702 N31701 N31702 10
D31702 N31702 0 diode
R31703 N31702 N31703 10
D31703 N31703 0 diode
R31704 N31703 N31704 10
D31704 N31704 0 diode
R31705 N31704 N31705 10
D31705 N31705 0 diode
R31706 N31705 N31706 10
D31706 N31706 0 diode
R31707 N31706 N31707 10
D31707 N31707 0 diode
R31708 N31707 N31708 10
D31708 N31708 0 diode
R31709 N31708 N31709 10
D31709 N31709 0 diode
R31710 N31709 N31710 10
D31710 N31710 0 diode
R31711 N31710 N31711 10
D31711 N31711 0 diode
R31712 N31711 N31712 10
D31712 N31712 0 diode
R31713 N31712 N31713 10
D31713 N31713 0 diode
R31714 N31713 N31714 10
D31714 N31714 0 diode
R31715 N31714 N31715 10
D31715 N31715 0 diode
R31716 N31715 N31716 10
D31716 N31716 0 diode
R31717 N31716 N31717 10
D31717 N31717 0 diode
R31718 N31717 N31718 10
D31718 N31718 0 diode
R31719 N31718 N31719 10
D31719 N31719 0 diode
R31720 N31719 N31720 10
D31720 N31720 0 diode
R31721 N31720 N31721 10
D31721 N31721 0 diode
R31722 N31721 N31722 10
D31722 N31722 0 diode
R31723 N31722 N31723 10
D31723 N31723 0 diode
R31724 N31723 N31724 10
D31724 N31724 0 diode
R31725 N31724 N31725 10
D31725 N31725 0 diode
R31726 N31725 N31726 10
D31726 N31726 0 diode
R31727 N31726 N31727 10
D31727 N31727 0 diode
R31728 N31727 N31728 10
D31728 N31728 0 diode
R31729 N31728 N31729 10
D31729 N31729 0 diode
R31730 N31729 N31730 10
D31730 N31730 0 diode
R31731 N31730 N31731 10
D31731 N31731 0 diode
R31732 N31731 N31732 10
D31732 N31732 0 diode
R31733 N31732 N31733 10
D31733 N31733 0 diode
R31734 N31733 N31734 10
D31734 N31734 0 diode
R31735 N31734 N31735 10
D31735 N31735 0 diode
R31736 N31735 N31736 10
D31736 N31736 0 diode
R31737 N31736 N31737 10
D31737 N31737 0 diode
R31738 N31737 N31738 10
D31738 N31738 0 diode
R31739 N31738 N31739 10
D31739 N31739 0 diode
R31740 N31739 N31740 10
D31740 N31740 0 diode
R31741 N31740 N31741 10
D31741 N31741 0 diode
R31742 N31741 N31742 10
D31742 N31742 0 diode
R31743 N31742 N31743 10
D31743 N31743 0 diode
R31744 N31743 N31744 10
D31744 N31744 0 diode
R31745 N31744 N31745 10
D31745 N31745 0 diode
R31746 N31745 N31746 10
D31746 N31746 0 diode
R31747 N31746 N31747 10
D31747 N31747 0 diode
R31748 N31747 N31748 10
D31748 N31748 0 diode
R31749 N31748 N31749 10
D31749 N31749 0 diode
R31750 N31749 N31750 10
D31750 N31750 0 diode
R31751 N31750 N31751 10
D31751 N31751 0 diode
R31752 N31751 N31752 10
D31752 N31752 0 diode
R31753 N31752 N31753 10
D31753 N31753 0 diode
R31754 N31753 N31754 10
D31754 N31754 0 diode
R31755 N31754 N31755 10
D31755 N31755 0 diode
R31756 N31755 N31756 10
D31756 N31756 0 diode
R31757 N31756 N31757 10
D31757 N31757 0 diode
R31758 N31757 N31758 10
D31758 N31758 0 diode
R31759 N31758 N31759 10
D31759 N31759 0 diode
R31760 N31759 N31760 10
D31760 N31760 0 diode
R31761 N31760 N31761 10
D31761 N31761 0 diode
R31762 N31761 N31762 10
D31762 N31762 0 diode
R31763 N31762 N31763 10
D31763 N31763 0 diode
R31764 N31763 N31764 10
D31764 N31764 0 diode
R31765 N31764 N31765 10
D31765 N31765 0 diode
R31766 N31765 N31766 10
D31766 N31766 0 diode
R31767 N31766 N31767 10
D31767 N31767 0 diode
R31768 N31767 N31768 10
D31768 N31768 0 diode
R31769 N31768 N31769 10
D31769 N31769 0 diode
R31770 N31769 N31770 10
D31770 N31770 0 diode
R31771 N31770 N31771 10
D31771 N31771 0 diode
R31772 N31771 N31772 10
D31772 N31772 0 diode
R31773 N31772 N31773 10
D31773 N31773 0 diode
R31774 N31773 N31774 10
D31774 N31774 0 diode
R31775 N31774 N31775 10
D31775 N31775 0 diode
R31776 N31775 N31776 10
D31776 N31776 0 diode
R31777 N31776 N31777 10
D31777 N31777 0 diode
R31778 N31777 N31778 10
D31778 N31778 0 diode
R31779 N31778 N31779 10
D31779 N31779 0 diode
R31780 N31779 N31780 10
D31780 N31780 0 diode
R31781 N31780 N31781 10
D31781 N31781 0 diode
R31782 N31781 N31782 10
D31782 N31782 0 diode
R31783 N31782 N31783 10
D31783 N31783 0 diode
R31784 N31783 N31784 10
D31784 N31784 0 diode
R31785 N31784 N31785 10
D31785 N31785 0 diode
R31786 N31785 N31786 10
D31786 N31786 0 diode
R31787 N31786 N31787 10
D31787 N31787 0 diode
R31788 N31787 N31788 10
D31788 N31788 0 diode
R31789 N31788 N31789 10
D31789 N31789 0 diode
R31790 N31789 N31790 10
D31790 N31790 0 diode
R31791 N31790 N31791 10
D31791 N31791 0 diode
R31792 N31791 N31792 10
D31792 N31792 0 diode
R31793 N31792 N31793 10
D31793 N31793 0 diode
R31794 N31793 N31794 10
D31794 N31794 0 diode
R31795 N31794 N31795 10
D31795 N31795 0 diode
R31796 N31795 N31796 10
D31796 N31796 0 diode
R31797 N31796 N31797 10
D31797 N31797 0 diode
R31798 N31797 N31798 10
D31798 N31798 0 diode
R31799 N31798 N31799 10
D31799 N31799 0 diode
R31800 N31799 N31800 10
D31800 N31800 0 diode
R31801 N31800 N31801 10
D31801 N31801 0 diode
R31802 N31801 N31802 10
D31802 N31802 0 diode
R31803 N31802 N31803 10
D31803 N31803 0 diode
R31804 N31803 N31804 10
D31804 N31804 0 diode
R31805 N31804 N31805 10
D31805 N31805 0 diode
R31806 N31805 N31806 10
D31806 N31806 0 diode
R31807 N31806 N31807 10
D31807 N31807 0 diode
R31808 N31807 N31808 10
D31808 N31808 0 diode
R31809 N31808 N31809 10
D31809 N31809 0 diode
R31810 N31809 N31810 10
D31810 N31810 0 diode
R31811 N31810 N31811 10
D31811 N31811 0 diode
R31812 N31811 N31812 10
D31812 N31812 0 diode
R31813 N31812 N31813 10
D31813 N31813 0 diode
R31814 N31813 N31814 10
D31814 N31814 0 diode
R31815 N31814 N31815 10
D31815 N31815 0 diode
R31816 N31815 N31816 10
D31816 N31816 0 diode
R31817 N31816 N31817 10
D31817 N31817 0 diode
R31818 N31817 N31818 10
D31818 N31818 0 diode
R31819 N31818 N31819 10
D31819 N31819 0 diode
R31820 N31819 N31820 10
D31820 N31820 0 diode
R31821 N31820 N31821 10
D31821 N31821 0 diode
R31822 N31821 N31822 10
D31822 N31822 0 diode
R31823 N31822 N31823 10
D31823 N31823 0 diode
R31824 N31823 N31824 10
D31824 N31824 0 diode
R31825 N31824 N31825 10
D31825 N31825 0 diode
R31826 N31825 N31826 10
D31826 N31826 0 diode
R31827 N31826 N31827 10
D31827 N31827 0 diode
R31828 N31827 N31828 10
D31828 N31828 0 diode
R31829 N31828 N31829 10
D31829 N31829 0 diode
R31830 N31829 N31830 10
D31830 N31830 0 diode
R31831 N31830 N31831 10
D31831 N31831 0 diode
R31832 N31831 N31832 10
D31832 N31832 0 diode
R31833 N31832 N31833 10
D31833 N31833 0 diode
R31834 N31833 N31834 10
D31834 N31834 0 diode
R31835 N31834 N31835 10
D31835 N31835 0 diode
R31836 N31835 N31836 10
D31836 N31836 0 diode
R31837 N31836 N31837 10
D31837 N31837 0 diode
R31838 N31837 N31838 10
D31838 N31838 0 diode
R31839 N31838 N31839 10
D31839 N31839 0 diode
R31840 N31839 N31840 10
D31840 N31840 0 diode
R31841 N31840 N31841 10
D31841 N31841 0 diode
R31842 N31841 N31842 10
D31842 N31842 0 diode
R31843 N31842 N31843 10
D31843 N31843 0 diode
R31844 N31843 N31844 10
D31844 N31844 0 diode
R31845 N31844 N31845 10
D31845 N31845 0 diode
R31846 N31845 N31846 10
D31846 N31846 0 diode
R31847 N31846 N31847 10
D31847 N31847 0 diode
R31848 N31847 N31848 10
D31848 N31848 0 diode
R31849 N31848 N31849 10
D31849 N31849 0 diode
R31850 N31849 N31850 10
D31850 N31850 0 diode
R31851 N31850 N31851 10
D31851 N31851 0 diode
R31852 N31851 N31852 10
D31852 N31852 0 diode
R31853 N31852 N31853 10
D31853 N31853 0 diode
R31854 N31853 N31854 10
D31854 N31854 0 diode
R31855 N31854 N31855 10
D31855 N31855 0 diode
R31856 N31855 N31856 10
D31856 N31856 0 diode
R31857 N31856 N31857 10
D31857 N31857 0 diode
R31858 N31857 N31858 10
D31858 N31858 0 diode
R31859 N31858 N31859 10
D31859 N31859 0 diode
R31860 N31859 N31860 10
D31860 N31860 0 diode
R31861 N31860 N31861 10
D31861 N31861 0 diode
R31862 N31861 N31862 10
D31862 N31862 0 diode
R31863 N31862 N31863 10
D31863 N31863 0 diode
R31864 N31863 N31864 10
D31864 N31864 0 diode
R31865 N31864 N31865 10
D31865 N31865 0 diode
R31866 N31865 N31866 10
D31866 N31866 0 diode
R31867 N31866 N31867 10
D31867 N31867 0 diode
R31868 N31867 N31868 10
D31868 N31868 0 diode
R31869 N31868 N31869 10
D31869 N31869 0 diode
R31870 N31869 N31870 10
D31870 N31870 0 diode
R31871 N31870 N31871 10
D31871 N31871 0 diode
R31872 N31871 N31872 10
D31872 N31872 0 diode
R31873 N31872 N31873 10
D31873 N31873 0 diode
R31874 N31873 N31874 10
D31874 N31874 0 diode
R31875 N31874 N31875 10
D31875 N31875 0 diode
R31876 N31875 N31876 10
D31876 N31876 0 diode
R31877 N31876 N31877 10
D31877 N31877 0 diode
R31878 N31877 N31878 10
D31878 N31878 0 diode
R31879 N31878 N31879 10
D31879 N31879 0 diode
R31880 N31879 N31880 10
D31880 N31880 0 diode
R31881 N31880 N31881 10
D31881 N31881 0 diode
R31882 N31881 N31882 10
D31882 N31882 0 diode
R31883 N31882 N31883 10
D31883 N31883 0 diode
R31884 N31883 N31884 10
D31884 N31884 0 diode
R31885 N31884 N31885 10
D31885 N31885 0 diode
R31886 N31885 N31886 10
D31886 N31886 0 diode
R31887 N31886 N31887 10
D31887 N31887 0 diode
R31888 N31887 N31888 10
D31888 N31888 0 diode
R31889 N31888 N31889 10
D31889 N31889 0 diode
R31890 N31889 N31890 10
D31890 N31890 0 diode
R31891 N31890 N31891 10
D31891 N31891 0 diode
R31892 N31891 N31892 10
D31892 N31892 0 diode
R31893 N31892 N31893 10
D31893 N31893 0 diode
R31894 N31893 N31894 10
D31894 N31894 0 diode
R31895 N31894 N31895 10
D31895 N31895 0 diode
R31896 N31895 N31896 10
D31896 N31896 0 diode
R31897 N31896 N31897 10
D31897 N31897 0 diode
R31898 N31897 N31898 10
D31898 N31898 0 diode
R31899 N31898 N31899 10
D31899 N31899 0 diode
R31900 N31899 N31900 10
D31900 N31900 0 diode
R31901 N31900 N31901 10
D31901 N31901 0 diode
R31902 N31901 N31902 10
D31902 N31902 0 diode
R31903 N31902 N31903 10
D31903 N31903 0 diode
R31904 N31903 N31904 10
D31904 N31904 0 diode
R31905 N31904 N31905 10
D31905 N31905 0 diode
R31906 N31905 N31906 10
D31906 N31906 0 diode
R31907 N31906 N31907 10
D31907 N31907 0 diode
R31908 N31907 N31908 10
D31908 N31908 0 diode
R31909 N31908 N31909 10
D31909 N31909 0 diode
R31910 N31909 N31910 10
D31910 N31910 0 diode
R31911 N31910 N31911 10
D31911 N31911 0 diode
R31912 N31911 N31912 10
D31912 N31912 0 diode
R31913 N31912 N31913 10
D31913 N31913 0 diode
R31914 N31913 N31914 10
D31914 N31914 0 diode
R31915 N31914 N31915 10
D31915 N31915 0 diode
R31916 N31915 N31916 10
D31916 N31916 0 diode
R31917 N31916 N31917 10
D31917 N31917 0 diode
R31918 N31917 N31918 10
D31918 N31918 0 diode
R31919 N31918 N31919 10
D31919 N31919 0 diode
R31920 N31919 N31920 10
D31920 N31920 0 diode
R31921 N31920 N31921 10
D31921 N31921 0 diode
R31922 N31921 N31922 10
D31922 N31922 0 diode
R31923 N31922 N31923 10
D31923 N31923 0 diode
R31924 N31923 N31924 10
D31924 N31924 0 diode
R31925 N31924 N31925 10
D31925 N31925 0 diode
R31926 N31925 N31926 10
D31926 N31926 0 diode
R31927 N31926 N31927 10
D31927 N31927 0 diode
R31928 N31927 N31928 10
D31928 N31928 0 diode
R31929 N31928 N31929 10
D31929 N31929 0 diode
R31930 N31929 N31930 10
D31930 N31930 0 diode
R31931 N31930 N31931 10
D31931 N31931 0 diode
R31932 N31931 N31932 10
D31932 N31932 0 diode
R31933 N31932 N31933 10
D31933 N31933 0 diode
R31934 N31933 N31934 10
D31934 N31934 0 diode
R31935 N31934 N31935 10
D31935 N31935 0 diode
R31936 N31935 N31936 10
D31936 N31936 0 diode
R31937 N31936 N31937 10
D31937 N31937 0 diode
R31938 N31937 N31938 10
D31938 N31938 0 diode
R31939 N31938 N31939 10
D31939 N31939 0 diode
R31940 N31939 N31940 10
D31940 N31940 0 diode
R31941 N31940 N31941 10
D31941 N31941 0 diode
R31942 N31941 N31942 10
D31942 N31942 0 diode
R31943 N31942 N31943 10
D31943 N31943 0 diode
R31944 N31943 N31944 10
D31944 N31944 0 diode
R31945 N31944 N31945 10
D31945 N31945 0 diode
R31946 N31945 N31946 10
D31946 N31946 0 diode
R31947 N31946 N31947 10
D31947 N31947 0 diode
R31948 N31947 N31948 10
D31948 N31948 0 diode
R31949 N31948 N31949 10
D31949 N31949 0 diode
R31950 N31949 N31950 10
D31950 N31950 0 diode
R31951 N31950 N31951 10
D31951 N31951 0 diode
R31952 N31951 N31952 10
D31952 N31952 0 diode
R31953 N31952 N31953 10
D31953 N31953 0 diode
R31954 N31953 N31954 10
D31954 N31954 0 diode
R31955 N31954 N31955 10
D31955 N31955 0 diode
R31956 N31955 N31956 10
D31956 N31956 0 diode
R31957 N31956 N31957 10
D31957 N31957 0 diode
R31958 N31957 N31958 10
D31958 N31958 0 diode
R31959 N31958 N31959 10
D31959 N31959 0 diode
R31960 N31959 N31960 10
D31960 N31960 0 diode
R31961 N31960 N31961 10
D31961 N31961 0 diode
R31962 N31961 N31962 10
D31962 N31962 0 diode
R31963 N31962 N31963 10
D31963 N31963 0 diode
R31964 N31963 N31964 10
D31964 N31964 0 diode
R31965 N31964 N31965 10
D31965 N31965 0 diode
R31966 N31965 N31966 10
D31966 N31966 0 diode
R31967 N31966 N31967 10
D31967 N31967 0 diode
R31968 N31967 N31968 10
D31968 N31968 0 diode
R31969 N31968 N31969 10
D31969 N31969 0 diode
R31970 N31969 N31970 10
D31970 N31970 0 diode
R31971 N31970 N31971 10
D31971 N31971 0 diode
R31972 N31971 N31972 10
D31972 N31972 0 diode
R31973 N31972 N31973 10
D31973 N31973 0 diode
R31974 N31973 N31974 10
D31974 N31974 0 diode
R31975 N31974 N31975 10
D31975 N31975 0 diode
R31976 N31975 N31976 10
D31976 N31976 0 diode
R31977 N31976 N31977 10
D31977 N31977 0 diode
R31978 N31977 N31978 10
D31978 N31978 0 diode
R31979 N31978 N31979 10
D31979 N31979 0 diode
R31980 N31979 N31980 10
D31980 N31980 0 diode
R31981 N31980 N31981 10
D31981 N31981 0 diode
R31982 N31981 N31982 10
D31982 N31982 0 diode
R31983 N31982 N31983 10
D31983 N31983 0 diode
R31984 N31983 N31984 10
D31984 N31984 0 diode
R31985 N31984 N31985 10
D31985 N31985 0 diode
R31986 N31985 N31986 10
D31986 N31986 0 diode
R31987 N31986 N31987 10
D31987 N31987 0 diode
R31988 N31987 N31988 10
D31988 N31988 0 diode
R31989 N31988 N31989 10
D31989 N31989 0 diode
R31990 N31989 N31990 10
D31990 N31990 0 diode
R31991 N31990 N31991 10
D31991 N31991 0 diode
R31992 N31991 N31992 10
D31992 N31992 0 diode
R31993 N31992 N31993 10
D31993 N31993 0 diode
R31994 N31993 N31994 10
D31994 N31994 0 diode
R31995 N31994 N31995 10
D31995 N31995 0 diode
R31996 N31995 N31996 10
D31996 N31996 0 diode
R31997 N31996 N31997 10
D31997 N31997 0 diode
R31998 N31997 N31998 10
D31998 N31998 0 diode
R31999 N31998 N31999 10
D31999 N31999 0 diode
R32000 N31999 N32000 10
D32000 N32000 0 diode
R32001 N32000 N32001 10
D32001 N32001 0 diode
R32002 N32001 N32002 10
D32002 N32002 0 diode
R32003 N32002 N32003 10
D32003 N32003 0 diode
R32004 N32003 N32004 10
D32004 N32004 0 diode
R32005 N32004 N32005 10
D32005 N32005 0 diode
R32006 N32005 N32006 10
D32006 N32006 0 diode
R32007 N32006 N32007 10
D32007 N32007 0 diode
R32008 N32007 N32008 10
D32008 N32008 0 diode
R32009 N32008 N32009 10
D32009 N32009 0 diode
R32010 N32009 N32010 10
D32010 N32010 0 diode
R32011 N32010 N32011 10
D32011 N32011 0 diode
R32012 N32011 N32012 10
D32012 N32012 0 diode
R32013 N32012 N32013 10
D32013 N32013 0 diode
R32014 N32013 N32014 10
D32014 N32014 0 diode
R32015 N32014 N32015 10
D32015 N32015 0 diode
R32016 N32015 N32016 10
D32016 N32016 0 diode
R32017 N32016 N32017 10
D32017 N32017 0 diode
R32018 N32017 N32018 10
D32018 N32018 0 diode
R32019 N32018 N32019 10
D32019 N32019 0 diode
R32020 N32019 N32020 10
D32020 N32020 0 diode
R32021 N32020 N32021 10
D32021 N32021 0 diode
R32022 N32021 N32022 10
D32022 N32022 0 diode
R32023 N32022 N32023 10
D32023 N32023 0 diode
R32024 N32023 N32024 10
D32024 N32024 0 diode
R32025 N32024 N32025 10
D32025 N32025 0 diode
R32026 N32025 N32026 10
D32026 N32026 0 diode
R32027 N32026 N32027 10
D32027 N32027 0 diode
R32028 N32027 N32028 10
D32028 N32028 0 diode
R32029 N32028 N32029 10
D32029 N32029 0 diode
R32030 N32029 N32030 10
D32030 N32030 0 diode
R32031 N32030 N32031 10
D32031 N32031 0 diode
R32032 N32031 N32032 10
D32032 N32032 0 diode
R32033 N32032 N32033 10
D32033 N32033 0 diode
R32034 N32033 N32034 10
D32034 N32034 0 diode
R32035 N32034 N32035 10
D32035 N32035 0 diode
R32036 N32035 N32036 10
D32036 N32036 0 diode
R32037 N32036 N32037 10
D32037 N32037 0 diode
R32038 N32037 N32038 10
D32038 N32038 0 diode
R32039 N32038 N32039 10
D32039 N32039 0 diode
R32040 N32039 N32040 10
D32040 N32040 0 diode
R32041 N32040 N32041 10
D32041 N32041 0 diode
R32042 N32041 N32042 10
D32042 N32042 0 diode
R32043 N32042 N32043 10
D32043 N32043 0 diode
R32044 N32043 N32044 10
D32044 N32044 0 diode
R32045 N32044 N32045 10
D32045 N32045 0 diode
R32046 N32045 N32046 10
D32046 N32046 0 diode
R32047 N32046 N32047 10
D32047 N32047 0 diode
R32048 N32047 N32048 10
D32048 N32048 0 diode
R32049 N32048 N32049 10
D32049 N32049 0 diode
R32050 N32049 N32050 10
D32050 N32050 0 diode
R32051 N32050 N32051 10
D32051 N32051 0 diode
R32052 N32051 N32052 10
D32052 N32052 0 diode
R32053 N32052 N32053 10
D32053 N32053 0 diode
R32054 N32053 N32054 10
D32054 N32054 0 diode
R32055 N32054 N32055 10
D32055 N32055 0 diode
R32056 N32055 N32056 10
D32056 N32056 0 diode
R32057 N32056 N32057 10
D32057 N32057 0 diode
R32058 N32057 N32058 10
D32058 N32058 0 diode
R32059 N32058 N32059 10
D32059 N32059 0 diode
R32060 N32059 N32060 10
D32060 N32060 0 diode
R32061 N32060 N32061 10
D32061 N32061 0 diode
R32062 N32061 N32062 10
D32062 N32062 0 diode
R32063 N32062 N32063 10
D32063 N32063 0 diode
R32064 N32063 N32064 10
D32064 N32064 0 diode
R32065 N32064 N32065 10
D32065 N32065 0 diode
R32066 N32065 N32066 10
D32066 N32066 0 diode
R32067 N32066 N32067 10
D32067 N32067 0 diode
R32068 N32067 N32068 10
D32068 N32068 0 diode
R32069 N32068 N32069 10
D32069 N32069 0 diode
R32070 N32069 N32070 10
D32070 N32070 0 diode
R32071 N32070 N32071 10
D32071 N32071 0 diode
R32072 N32071 N32072 10
D32072 N32072 0 diode
R32073 N32072 N32073 10
D32073 N32073 0 diode
R32074 N32073 N32074 10
D32074 N32074 0 diode
R32075 N32074 N32075 10
D32075 N32075 0 diode
R32076 N32075 N32076 10
D32076 N32076 0 diode
R32077 N32076 N32077 10
D32077 N32077 0 diode
R32078 N32077 N32078 10
D32078 N32078 0 diode
R32079 N32078 N32079 10
D32079 N32079 0 diode
R32080 N32079 N32080 10
D32080 N32080 0 diode
R32081 N32080 N32081 10
D32081 N32081 0 diode
R32082 N32081 N32082 10
D32082 N32082 0 diode
R32083 N32082 N32083 10
D32083 N32083 0 diode
R32084 N32083 N32084 10
D32084 N32084 0 diode
R32085 N32084 N32085 10
D32085 N32085 0 diode
R32086 N32085 N32086 10
D32086 N32086 0 diode
R32087 N32086 N32087 10
D32087 N32087 0 diode
R32088 N32087 N32088 10
D32088 N32088 0 diode
R32089 N32088 N32089 10
D32089 N32089 0 diode
R32090 N32089 N32090 10
D32090 N32090 0 diode
R32091 N32090 N32091 10
D32091 N32091 0 diode
R32092 N32091 N32092 10
D32092 N32092 0 diode
R32093 N32092 N32093 10
D32093 N32093 0 diode
R32094 N32093 N32094 10
D32094 N32094 0 diode
R32095 N32094 N32095 10
D32095 N32095 0 diode
R32096 N32095 N32096 10
D32096 N32096 0 diode
R32097 N32096 N32097 10
D32097 N32097 0 diode
R32098 N32097 N32098 10
D32098 N32098 0 diode
R32099 N32098 N32099 10
D32099 N32099 0 diode
R32100 N32099 N32100 10
D32100 N32100 0 diode
R32101 N32100 N32101 10
D32101 N32101 0 diode
R32102 N32101 N32102 10
D32102 N32102 0 diode
R32103 N32102 N32103 10
D32103 N32103 0 diode
R32104 N32103 N32104 10
D32104 N32104 0 diode
R32105 N32104 N32105 10
D32105 N32105 0 diode
R32106 N32105 N32106 10
D32106 N32106 0 diode
R32107 N32106 N32107 10
D32107 N32107 0 diode
R32108 N32107 N32108 10
D32108 N32108 0 diode
R32109 N32108 N32109 10
D32109 N32109 0 diode
R32110 N32109 N32110 10
D32110 N32110 0 diode
R32111 N32110 N32111 10
D32111 N32111 0 diode
R32112 N32111 N32112 10
D32112 N32112 0 diode
R32113 N32112 N32113 10
D32113 N32113 0 diode
R32114 N32113 N32114 10
D32114 N32114 0 diode
R32115 N32114 N32115 10
D32115 N32115 0 diode
R32116 N32115 N32116 10
D32116 N32116 0 diode
R32117 N32116 N32117 10
D32117 N32117 0 diode
R32118 N32117 N32118 10
D32118 N32118 0 diode
R32119 N32118 N32119 10
D32119 N32119 0 diode
R32120 N32119 N32120 10
D32120 N32120 0 diode
R32121 N32120 N32121 10
D32121 N32121 0 diode
R32122 N32121 N32122 10
D32122 N32122 0 diode
R32123 N32122 N32123 10
D32123 N32123 0 diode
R32124 N32123 N32124 10
D32124 N32124 0 diode
R32125 N32124 N32125 10
D32125 N32125 0 diode
R32126 N32125 N32126 10
D32126 N32126 0 diode
R32127 N32126 N32127 10
D32127 N32127 0 diode
R32128 N32127 N32128 10
D32128 N32128 0 diode
R32129 N32128 N32129 10
D32129 N32129 0 diode
R32130 N32129 N32130 10
D32130 N32130 0 diode
R32131 N32130 N32131 10
D32131 N32131 0 diode
R32132 N32131 N32132 10
D32132 N32132 0 diode
R32133 N32132 N32133 10
D32133 N32133 0 diode
R32134 N32133 N32134 10
D32134 N32134 0 diode
R32135 N32134 N32135 10
D32135 N32135 0 diode
R32136 N32135 N32136 10
D32136 N32136 0 diode
R32137 N32136 N32137 10
D32137 N32137 0 diode
R32138 N32137 N32138 10
D32138 N32138 0 diode
R32139 N32138 N32139 10
D32139 N32139 0 diode
R32140 N32139 N32140 10
D32140 N32140 0 diode
R32141 N32140 N32141 10
D32141 N32141 0 diode
R32142 N32141 N32142 10
D32142 N32142 0 diode
R32143 N32142 N32143 10
D32143 N32143 0 diode
R32144 N32143 N32144 10
D32144 N32144 0 diode
R32145 N32144 N32145 10
D32145 N32145 0 diode
R32146 N32145 N32146 10
D32146 N32146 0 diode
R32147 N32146 N32147 10
D32147 N32147 0 diode
R32148 N32147 N32148 10
D32148 N32148 0 diode
R32149 N32148 N32149 10
D32149 N32149 0 diode
R32150 N32149 N32150 10
D32150 N32150 0 diode
R32151 N32150 N32151 10
D32151 N32151 0 diode
R32152 N32151 N32152 10
D32152 N32152 0 diode
R32153 N32152 N32153 10
D32153 N32153 0 diode
R32154 N32153 N32154 10
D32154 N32154 0 diode
R32155 N32154 N32155 10
D32155 N32155 0 diode
R32156 N32155 N32156 10
D32156 N32156 0 diode
R32157 N32156 N32157 10
D32157 N32157 0 diode
R32158 N32157 N32158 10
D32158 N32158 0 diode
R32159 N32158 N32159 10
D32159 N32159 0 diode
R32160 N32159 N32160 10
D32160 N32160 0 diode
R32161 N32160 N32161 10
D32161 N32161 0 diode
R32162 N32161 N32162 10
D32162 N32162 0 diode
R32163 N32162 N32163 10
D32163 N32163 0 diode
R32164 N32163 N32164 10
D32164 N32164 0 diode
R32165 N32164 N32165 10
D32165 N32165 0 diode
R32166 N32165 N32166 10
D32166 N32166 0 diode
R32167 N32166 N32167 10
D32167 N32167 0 diode
R32168 N32167 N32168 10
D32168 N32168 0 diode
R32169 N32168 N32169 10
D32169 N32169 0 diode
R32170 N32169 N32170 10
D32170 N32170 0 diode
R32171 N32170 N32171 10
D32171 N32171 0 diode
R32172 N32171 N32172 10
D32172 N32172 0 diode
R32173 N32172 N32173 10
D32173 N32173 0 diode
R32174 N32173 N32174 10
D32174 N32174 0 diode
R32175 N32174 N32175 10
D32175 N32175 0 diode
R32176 N32175 N32176 10
D32176 N32176 0 diode
R32177 N32176 N32177 10
D32177 N32177 0 diode
R32178 N32177 N32178 10
D32178 N32178 0 diode
R32179 N32178 N32179 10
D32179 N32179 0 diode
R32180 N32179 N32180 10
D32180 N32180 0 diode
R32181 N32180 N32181 10
D32181 N32181 0 diode
R32182 N32181 N32182 10
D32182 N32182 0 diode
R32183 N32182 N32183 10
D32183 N32183 0 diode
R32184 N32183 N32184 10
D32184 N32184 0 diode
R32185 N32184 N32185 10
D32185 N32185 0 diode
R32186 N32185 N32186 10
D32186 N32186 0 diode
R32187 N32186 N32187 10
D32187 N32187 0 diode
R32188 N32187 N32188 10
D32188 N32188 0 diode
R32189 N32188 N32189 10
D32189 N32189 0 diode
R32190 N32189 N32190 10
D32190 N32190 0 diode
R32191 N32190 N32191 10
D32191 N32191 0 diode
R32192 N32191 N32192 10
D32192 N32192 0 diode
R32193 N32192 N32193 10
D32193 N32193 0 diode
R32194 N32193 N32194 10
D32194 N32194 0 diode
R32195 N32194 N32195 10
D32195 N32195 0 diode
R32196 N32195 N32196 10
D32196 N32196 0 diode
R32197 N32196 N32197 10
D32197 N32197 0 diode
R32198 N32197 N32198 10
D32198 N32198 0 diode
R32199 N32198 N32199 10
D32199 N32199 0 diode
R32200 N32199 N32200 10
D32200 N32200 0 diode
R32201 N32200 N32201 10
D32201 N32201 0 diode
R32202 N32201 N32202 10
D32202 N32202 0 diode
R32203 N32202 N32203 10
D32203 N32203 0 diode
R32204 N32203 N32204 10
D32204 N32204 0 diode
R32205 N32204 N32205 10
D32205 N32205 0 diode
R32206 N32205 N32206 10
D32206 N32206 0 diode
R32207 N32206 N32207 10
D32207 N32207 0 diode
R32208 N32207 N32208 10
D32208 N32208 0 diode
R32209 N32208 N32209 10
D32209 N32209 0 diode
R32210 N32209 N32210 10
D32210 N32210 0 diode
R32211 N32210 N32211 10
D32211 N32211 0 diode
R32212 N32211 N32212 10
D32212 N32212 0 diode
R32213 N32212 N32213 10
D32213 N32213 0 diode
R32214 N32213 N32214 10
D32214 N32214 0 diode
R32215 N32214 N32215 10
D32215 N32215 0 diode
R32216 N32215 N32216 10
D32216 N32216 0 diode
R32217 N32216 N32217 10
D32217 N32217 0 diode
R32218 N32217 N32218 10
D32218 N32218 0 diode
R32219 N32218 N32219 10
D32219 N32219 0 diode
R32220 N32219 N32220 10
D32220 N32220 0 diode
R32221 N32220 N32221 10
D32221 N32221 0 diode
R32222 N32221 N32222 10
D32222 N32222 0 diode
R32223 N32222 N32223 10
D32223 N32223 0 diode
R32224 N32223 N32224 10
D32224 N32224 0 diode
R32225 N32224 N32225 10
D32225 N32225 0 diode
R32226 N32225 N32226 10
D32226 N32226 0 diode
R32227 N32226 N32227 10
D32227 N32227 0 diode
R32228 N32227 N32228 10
D32228 N32228 0 diode
R32229 N32228 N32229 10
D32229 N32229 0 diode
R32230 N32229 N32230 10
D32230 N32230 0 diode
R32231 N32230 N32231 10
D32231 N32231 0 diode
R32232 N32231 N32232 10
D32232 N32232 0 diode
R32233 N32232 N32233 10
D32233 N32233 0 diode
R32234 N32233 N32234 10
D32234 N32234 0 diode
R32235 N32234 N32235 10
D32235 N32235 0 diode
R32236 N32235 N32236 10
D32236 N32236 0 diode
R32237 N32236 N32237 10
D32237 N32237 0 diode
R32238 N32237 N32238 10
D32238 N32238 0 diode
R32239 N32238 N32239 10
D32239 N32239 0 diode
R32240 N32239 N32240 10
D32240 N32240 0 diode
R32241 N32240 N32241 10
D32241 N32241 0 diode
R32242 N32241 N32242 10
D32242 N32242 0 diode
R32243 N32242 N32243 10
D32243 N32243 0 diode
R32244 N32243 N32244 10
D32244 N32244 0 diode
R32245 N32244 N32245 10
D32245 N32245 0 diode
R32246 N32245 N32246 10
D32246 N32246 0 diode
R32247 N32246 N32247 10
D32247 N32247 0 diode
R32248 N32247 N32248 10
D32248 N32248 0 diode
R32249 N32248 N32249 10
D32249 N32249 0 diode
R32250 N32249 N32250 10
D32250 N32250 0 diode
R32251 N32250 N32251 10
D32251 N32251 0 diode
R32252 N32251 N32252 10
D32252 N32252 0 diode
R32253 N32252 N32253 10
D32253 N32253 0 diode
R32254 N32253 N32254 10
D32254 N32254 0 diode
R32255 N32254 N32255 10
D32255 N32255 0 diode
R32256 N32255 N32256 10
D32256 N32256 0 diode
R32257 N32256 N32257 10
D32257 N32257 0 diode
R32258 N32257 N32258 10
D32258 N32258 0 diode
R32259 N32258 N32259 10
D32259 N32259 0 diode
R32260 N32259 N32260 10
D32260 N32260 0 diode
R32261 N32260 N32261 10
D32261 N32261 0 diode
R32262 N32261 N32262 10
D32262 N32262 0 diode
R32263 N32262 N32263 10
D32263 N32263 0 diode
R32264 N32263 N32264 10
D32264 N32264 0 diode
R32265 N32264 N32265 10
D32265 N32265 0 diode
R32266 N32265 N32266 10
D32266 N32266 0 diode
R32267 N32266 N32267 10
D32267 N32267 0 diode
R32268 N32267 N32268 10
D32268 N32268 0 diode
R32269 N32268 N32269 10
D32269 N32269 0 diode
R32270 N32269 N32270 10
D32270 N32270 0 diode
R32271 N32270 N32271 10
D32271 N32271 0 diode
R32272 N32271 N32272 10
D32272 N32272 0 diode
R32273 N32272 N32273 10
D32273 N32273 0 diode
R32274 N32273 N32274 10
D32274 N32274 0 diode
R32275 N32274 N32275 10
D32275 N32275 0 diode
R32276 N32275 N32276 10
D32276 N32276 0 diode
R32277 N32276 N32277 10
D32277 N32277 0 diode
R32278 N32277 N32278 10
D32278 N32278 0 diode
R32279 N32278 N32279 10
D32279 N32279 0 diode
R32280 N32279 N32280 10
D32280 N32280 0 diode
R32281 N32280 N32281 10
D32281 N32281 0 diode
R32282 N32281 N32282 10
D32282 N32282 0 diode
R32283 N32282 N32283 10
D32283 N32283 0 diode
R32284 N32283 N32284 10
D32284 N32284 0 diode
R32285 N32284 N32285 10
D32285 N32285 0 diode
R32286 N32285 N32286 10
D32286 N32286 0 diode
R32287 N32286 N32287 10
D32287 N32287 0 diode
R32288 N32287 N32288 10
D32288 N32288 0 diode
R32289 N32288 N32289 10
D32289 N32289 0 diode
R32290 N32289 N32290 10
D32290 N32290 0 diode
R32291 N32290 N32291 10
D32291 N32291 0 diode
R32292 N32291 N32292 10
D32292 N32292 0 diode
R32293 N32292 N32293 10
D32293 N32293 0 diode
R32294 N32293 N32294 10
D32294 N32294 0 diode
R32295 N32294 N32295 10
D32295 N32295 0 diode
R32296 N32295 N32296 10
D32296 N32296 0 diode
R32297 N32296 N32297 10
D32297 N32297 0 diode
R32298 N32297 N32298 10
D32298 N32298 0 diode
R32299 N32298 N32299 10
D32299 N32299 0 diode
R32300 N32299 N32300 10
D32300 N32300 0 diode
R32301 N32300 N32301 10
D32301 N32301 0 diode
R32302 N32301 N32302 10
D32302 N32302 0 diode
R32303 N32302 N32303 10
D32303 N32303 0 diode
R32304 N32303 N32304 10
D32304 N32304 0 diode
R32305 N32304 N32305 10
D32305 N32305 0 diode
R32306 N32305 N32306 10
D32306 N32306 0 diode
R32307 N32306 N32307 10
D32307 N32307 0 diode
R32308 N32307 N32308 10
D32308 N32308 0 diode
R32309 N32308 N32309 10
D32309 N32309 0 diode
R32310 N32309 N32310 10
D32310 N32310 0 diode
R32311 N32310 N32311 10
D32311 N32311 0 diode
R32312 N32311 N32312 10
D32312 N32312 0 diode
R32313 N32312 N32313 10
D32313 N32313 0 diode
R32314 N32313 N32314 10
D32314 N32314 0 diode
R32315 N32314 N32315 10
D32315 N32315 0 diode
R32316 N32315 N32316 10
D32316 N32316 0 diode
R32317 N32316 N32317 10
D32317 N32317 0 diode
R32318 N32317 N32318 10
D32318 N32318 0 diode
R32319 N32318 N32319 10
D32319 N32319 0 diode
R32320 N32319 N32320 10
D32320 N32320 0 diode
R32321 N32320 N32321 10
D32321 N32321 0 diode
R32322 N32321 N32322 10
D32322 N32322 0 diode
R32323 N32322 N32323 10
D32323 N32323 0 diode
R32324 N32323 N32324 10
D32324 N32324 0 diode
R32325 N32324 N32325 10
D32325 N32325 0 diode
R32326 N32325 N32326 10
D32326 N32326 0 diode
R32327 N32326 N32327 10
D32327 N32327 0 diode
R32328 N32327 N32328 10
D32328 N32328 0 diode
R32329 N32328 N32329 10
D32329 N32329 0 diode
R32330 N32329 N32330 10
D32330 N32330 0 diode
R32331 N32330 N32331 10
D32331 N32331 0 diode
R32332 N32331 N32332 10
D32332 N32332 0 diode
R32333 N32332 N32333 10
D32333 N32333 0 diode
R32334 N32333 N32334 10
D32334 N32334 0 diode
R32335 N32334 N32335 10
D32335 N32335 0 diode
R32336 N32335 N32336 10
D32336 N32336 0 diode
R32337 N32336 N32337 10
D32337 N32337 0 diode
R32338 N32337 N32338 10
D32338 N32338 0 diode
R32339 N32338 N32339 10
D32339 N32339 0 diode
R32340 N32339 N32340 10
D32340 N32340 0 diode
R32341 N32340 N32341 10
D32341 N32341 0 diode
R32342 N32341 N32342 10
D32342 N32342 0 diode
R32343 N32342 N32343 10
D32343 N32343 0 diode
R32344 N32343 N32344 10
D32344 N32344 0 diode
R32345 N32344 N32345 10
D32345 N32345 0 diode
R32346 N32345 N32346 10
D32346 N32346 0 diode
R32347 N32346 N32347 10
D32347 N32347 0 diode
R32348 N32347 N32348 10
D32348 N32348 0 diode
R32349 N32348 N32349 10
D32349 N32349 0 diode
R32350 N32349 N32350 10
D32350 N32350 0 diode
R32351 N32350 N32351 10
D32351 N32351 0 diode
R32352 N32351 N32352 10
D32352 N32352 0 diode
R32353 N32352 N32353 10
D32353 N32353 0 diode
R32354 N32353 N32354 10
D32354 N32354 0 diode
R32355 N32354 N32355 10
D32355 N32355 0 diode
R32356 N32355 N32356 10
D32356 N32356 0 diode
R32357 N32356 N32357 10
D32357 N32357 0 diode
R32358 N32357 N32358 10
D32358 N32358 0 diode
R32359 N32358 N32359 10
D32359 N32359 0 diode
R32360 N32359 N32360 10
D32360 N32360 0 diode
R32361 N32360 N32361 10
D32361 N32361 0 diode
R32362 N32361 N32362 10
D32362 N32362 0 diode
R32363 N32362 N32363 10
D32363 N32363 0 diode
R32364 N32363 N32364 10
D32364 N32364 0 diode
R32365 N32364 N32365 10
D32365 N32365 0 diode
R32366 N32365 N32366 10
D32366 N32366 0 diode
R32367 N32366 N32367 10
D32367 N32367 0 diode
R32368 N32367 N32368 10
D32368 N32368 0 diode
R32369 N32368 N32369 10
D32369 N32369 0 diode
R32370 N32369 N32370 10
D32370 N32370 0 diode
R32371 N32370 N32371 10
D32371 N32371 0 diode
R32372 N32371 N32372 10
D32372 N32372 0 diode
R32373 N32372 N32373 10
D32373 N32373 0 diode
R32374 N32373 N32374 10
D32374 N32374 0 diode
R32375 N32374 N32375 10
D32375 N32375 0 diode
R32376 N32375 N32376 10
D32376 N32376 0 diode
R32377 N32376 N32377 10
D32377 N32377 0 diode
R32378 N32377 N32378 10
D32378 N32378 0 diode
R32379 N32378 N32379 10
D32379 N32379 0 diode
R32380 N32379 N32380 10
D32380 N32380 0 diode
R32381 N32380 N32381 10
D32381 N32381 0 diode
R32382 N32381 N32382 10
D32382 N32382 0 diode
R32383 N32382 N32383 10
D32383 N32383 0 diode
R32384 N32383 N32384 10
D32384 N32384 0 diode
R32385 N32384 N32385 10
D32385 N32385 0 diode
R32386 N32385 N32386 10
D32386 N32386 0 diode
R32387 N32386 N32387 10
D32387 N32387 0 diode
R32388 N32387 N32388 10
D32388 N32388 0 diode
R32389 N32388 N32389 10
D32389 N32389 0 diode
R32390 N32389 N32390 10
D32390 N32390 0 diode
R32391 N32390 N32391 10
D32391 N32391 0 diode
R32392 N32391 N32392 10
D32392 N32392 0 diode
R32393 N32392 N32393 10
D32393 N32393 0 diode
R32394 N32393 N32394 10
D32394 N32394 0 diode
R32395 N32394 N32395 10
D32395 N32395 0 diode
R32396 N32395 N32396 10
D32396 N32396 0 diode
R32397 N32396 N32397 10
D32397 N32397 0 diode
R32398 N32397 N32398 10
D32398 N32398 0 diode
R32399 N32398 N32399 10
D32399 N32399 0 diode
R32400 N32399 N32400 10
D32400 N32400 0 diode
R32401 N32400 N32401 10
D32401 N32401 0 diode
R32402 N32401 N32402 10
D32402 N32402 0 diode
R32403 N32402 N32403 10
D32403 N32403 0 diode
R32404 N32403 N32404 10
D32404 N32404 0 diode
R32405 N32404 N32405 10
D32405 N32405 0 diode
R32406 N32405 N32406 10
D32406 N32406 0 diode
R32407 N32406 N32407 10
D32407 N32407 0 diode
R32408 N32407 N32408 10
D32408 N32408 0 diode
R32409 N32408 N32409 10
D32409 N32409 0 diode
R32410 N32409 N32410 10
D32410 N32410 0 diode
R32411 N32410 N32411 10
D32411 N32411 0 diode
R32412 N32411 N32412 10
D32412 N32412 0 diode
R32413 N32412 N32413 10
D32413 N32413 0 diode
R32414 N32413 N32414 10
D32414 N32414 0 diode
R32415 N32414 N32415 10
D32415 N32415 0 diode
R32416 N32415 N32416 10
D32416 N32416 0 diode
R32417 N32416 N32417 10
D32417 N32417 0 diode
R32418 N32417 N32418 10
D32418 N32418 0 diode
R32419 N32418 N32419 10
D32419 N32419 0 diode
R32420 N32419 N32420 10
D32420 N32420 0 diode
R32421 N32420 N32421 10
D32421 N32421 0 diode
R32422 N32421 N32422 10
D32422 N32422 0 diode
R32423 N32422 N32423 10
D32423 N32423 0 diode
R32424 N32423 N32424 10
D32424 N32424 0 diode
R32425 N32424 N32425 10
D32425 N32425 0 diode
R32426 N32425 N32426 10
D32426 N32426 0 diode
R32427 N32426 N32427 10
D32427 N32427 0 diode
R32428 N32427 N32428 10
D32428 N32428 0 diode
R32429 N32428 N32429 10
D32429 N32429 0 diode
R32430 N32429 N32430 10
D32430 N32430 0 diode
R32431 N32430 N32431 10
D32431 N32431 0 diode
R32432 N32431 N32432 10
D32432 N32432 0 diode
R32433 N32432 N32433 10
D32433 N32433 0 diode
R32434 N32433 N32434 10
D32434 N32434 0 diode
R32435 N32434 N32435 10
D32435 N32435 0 diode
R32436 N32435 N32436 10
D32436 N32436 0 diode
R32437 N32436 N32437 10
D32437 N32437 0 diode
R32438 N32437 N32438 10
D32438 N32438 0 diode
R32439 N32438 N32439 10
D32439 N32439 0 diode
R32440 N32439 N32440 10
D32440 N32440 0 diode
R32441 N32440 N32441 10
D32441 N32441 0 diode
R32442 N32441 N32442 10
D32442 N32442 0 diode
R32443 N32442 N32443 10
D32443 N32443 0 diode
R32444 N32443 N32444 10
D32444 N32444 0 diode
R32445 N32444 N32445 10
D32445 N32445 0 diode
R32446 N32445 N32446 10
D32446 N32446 0 diode
R32447 N32446 N32447 10
D32447 N32447 0 diode
R32448 N32447 N32448 10
D32448 N32448 0 diode
R32449 N32448 N32449 10
D32449 N32449 0 diode
R32450 N32449 N32450 10
D32450 N32450 0 diode
R32451 N32450 N32451 10
D32451 N32451 0 diode
R32452 N32451 N32452 10
D32452 N32452 0 diode
R32453 N32452 N32453 10
D32453 N32453 0 diode
R32454 N32453 N32454 10
D32454 N32454 0 diode
R32455 N32454 N32455 10
D32455 N32455 0 diode
R32456 N32455 N32456 10
D32456 N32456 0 diode
R32457 N32456 N32457 10
D32457 N32457 0 diode
R32458 N32457 N32458 10
D32458 N32458 0 diode
R32459 N32458 N32459 10
D32459 N32459 0 diode
R32460 N32459 N32460 10
D32460 N32460 0 diode
R32461 N32460 N32461 10
D32461 N32461 0 diode
R32462 N32461 N32462 10
D32462 N32462 0 diode
R32463 N32462 N32463 10
D32463 N32463 0 diode
R32464 N32463 N32464 10
D32464 N32464 0 diode
R32465 N32464 N32465 10
D32465 N32465 0 diode
R32466 N32465 N32466 10
D32466 N32466 0 diode
R32467 N32466 N32467 10
D32467 N32467 0 diode
R32468 N32467 N32468 10
D32468 N32468 0 diode
R32469 N32468 N32469 10
D32469 N32469 0 diode
R32470 N32469 N32470 10
D32470 N32470 0 diode
R32471 N32470 N32471 10
D32471 N32471 0 diode
R32472 N32471 N32472 10
D32472 N32472 0 diode
R32473 N32472 N32473 10
D32473 N32473 0 diode
R32474 N32473 N32474 10
D32474 N32474 0 diode
R32475 N32474 N32475 10
D32475 N32475 0 diode
R32476 N32475 N32476 10
D32476 N32476 0 diode
R32477 N32476 N32477 10
D32477 N32477 0 diode
R32478 N32477 N32478 10
D32478 N32478 0 diode
R32479 N32478 N32479 10
D32479 N32479 0 diode
R32480 N32479 N32480 10
D32480 N32480 0 diode
R32481 N32480 N32481 10
D32481 N32481 0 diode
R32482 N32481 N32482 10
D32482 N32482 0 diode
R32483 N32482 N32483 10
D32483 N32483 0 diode
R32484 N32483 N32484 10
D32484 N32484 0 diode
R32485 N32484 N32485 10
D32485 N32485 0 diode
R32486 N32485 N32486 10
D32486 N32486 0 diode
R32487 N32486 N32487 10
D32487 N32487 0 diode
R32488 N32487 N32488 10
D32488 N32488 0 diode
R32489 N32488 N32489 10
D32489 N32489 0 diode
R32490 N32489 N32490 10
D32490 N32490 0 diode
R32491 N32490 N32491 10
D32491 N32491 0 diode
R32492 N32491 N32492 10
D32492 N32492 0 diode
R32493 N32492 N32493 10
D32493 N32493 0 diode
R32494 N32493 N32494 10
D32494 N32494 0 diode
R32495 N32494 N32495 10
D32495 N32495 0 diode
R32496 N32495 N32496 10
D32496 N32496 0 diode
R32497 N32496 N32497 10
D32497 N32497 0 diode
R32498 N32497 N32498 10
D32498 N32498 0 diode
R32499 N32498 N32499 10
D32499 N32499 0 diode
R32500 N32499 N32500 10
D32500 N32500 0 diode
R32501 N32500 N32501 10
D32501 N32501 0 diode
R32502 N32501 N32502 10
D32502 N32502 0 diode
R32503 N32502 N32503 10
D32503 N32503 0 diode
R32504 N32503 N32504 10
D32504 N32504 0 diode
R32505 N32504 N32505 10
D32505 N32505 0 diode
R32506 N32505 N32506 10
D32506 N32506 0 diode
R32507 N32506 N32507 10
D32507 N32507 0 diode
R32508 N32507 N32508 10
D32508 N32508 0 diode
R32509 N32508 N32509 10
D32509 N32509 0 diode
R32510 N32509 N32510 10
D32510 N32510 0 diode
R32511 N32510 N32511 10
D32511 N32511 0 diode
R32512 N32511 N32512 10
D32512 N32512 0 diode
R32513 N32512 N32513 10
D32513 N32513 0 diode
R32514 N32513 N32514 10
D32514 N32514 0 diode
R32515 N32514 N32515 10
D32515 N32515 0 diode
R32516 N32515 N32516 10
D32516 N32516 0 diode
R32517 N32516 N32517 10
D32517 N32517 0 diode
R32518 N32517 N32518 10
D32518 N32518 0 diode
R32519 N32518 N32519 10
D32519 N32519 0 diode
R32520 N32519 N32520 10
D32520 N32520 0 diode
R32521 N32520 N32521 10
D32521 N32521 0 diode
R32522 N32521 N32522 10
D32522 N32522 0 diode
R32523 N32522 N32523 10
D32523 N32523 0 diode
R32524 N32523 N32524 10
D32524 N32524 0 diode
R32525 N32524 N32525 10
D32525 N32525 0 diode
R32526 N32525 N32526 10
D32526 N32526 0 diode
R32527 N32526 N32527 10
D32527 N32527 0 diode
R32528 N32527 N32528 10
D32528 N32528 0 diode
R32529 N32528 N32529 10
D32529 N32529 0 diode
R32530 N32529 N32530 10
D32530 N32530 0 diode
R32531 N32530 N32531 10
D32531 N32531 0 diode
R32532 N32531 N32532 10
D32532 N32532 0 diode
R32533 N32532 N32533 10
D32533 N32533 0 diode
R32534 N32533 N32534 10
D32534 N32534 0 diode
R32535 N32534 N32535 10
D32535 N32535 0 diode
R32536 N32535 N32536 10
D32536 N32536 0 diode
R32537 N32536 N32537 10
D32537 N32537 0 diode
R32538 N32537 N32538 10
D32538 N32538 0 diode
R32539 N32538 N32539 10
D32539 N32539 0 diode
R32540 N32539 N32540 10
D32540 N32540 0 diode
R32541 N32540 N32541 10
D32541 N32541 0 diode
R32542 N32541 N32542 10
D32542 N32542 0 diode
R32543 N32542 N32543 10
D32543 N32543 0 diode
R32544 N32543 N32544 10
D32544 N32544 0 diode
R32545 N32544 N32545 10
D32545 N32545 0 diode
R32546 N32545 N32546 10
D32546 N32546 0 diode
R32547 N32546 N32547 10
D32547 N32547 0 diode
R32548 N32547 N32548 10
D32548 N32548 0 diode
R32549 N32548 N32549 10
D32549 N32549 0 diode
R32550 N32549 N32550 10
D32550 N32550 0 diode
R32551 N32550 N32551 10
D32551 N32551 0 diode
R32552 N32551 N32552 10
D32552 N32552 0 diode
R32553 N32552 N32553 10
D32553 N32553 0 diode
R32554 N32553 N32554 10
D32554 N32554 0 diode
R32555 N32554 N32555 10
D32555 N32555 0 diode
R32556 N32555 N32556 10
D32556 N32556 0 diode
R32557 N32556 N32557 10
D32557 N32557 0 diode
R32558 N32557 N32558 10
D32558 N32558 0 diode
R32559 N32558 N32559 10
D32559 N32559 0 diode
R32560 N32559 N32560 10
D32560 N32560 0 diode
R32561 N32560 N32561 10
D32561 N32561 0 diode
R32562 N32561 N32562 10
D32562 N32562 0 diode
R32563 N32562 N32563 10
D32563 N32563 0 diode
R32564 N32563 N32564 10
D32564 N32564 0 diode
R32565 N32564 N32565 10
D32565 N32565 0 diode
R32566 N32565 N32566 10
D32566 N32566 0 diode
R32567 N32566 N32567 10
D32567 N32567 0 diode
R32568 N32567 N32568 10
D32568 N32568 0 diode
R32569 N32568 N32569 10
D32569 N32569 0 diode
R32570 N32569 N32570 10
D32570 N32570 0 diode
R32571 N32570 N32571 10
D32571 N32571 0 diode
R32572 N32571 N32572 10
D32572 N32572 0 diode
R32573 N32572 N32573 10
D32573 N32573 0 diode
R32574 N32573 N32574 10
D32574 N32574 0 diode
R32575 N32574 N32575 10
D32575 N32575 0 diode
R32576 N32575 N32576 10
D32576 N32576 0 diode
R32577 N32576 N32577 10
D32577 N32577 0 diode
R32578 N32577 N32578 10
D32578 N32578 0 diode
R32579 N32578 N32579 10
D32579 N32579 0 diode
R32580 N32579 N32580 10
D32580 N32580 0 diode
R32581 N32580 N32581 10
D32581 N32581 0 diode
R32582 N32581 N32582 10
D32582 N32582 0 diode
R32583 N32582 N32583 10
D32583 N32583 0 diode
R32584 N32583 N32584 10
D32584 N32584 0 diode
R32585 N32584 N32585 10
D32585 N32585 0 diode
R32586 N32585 N32586 10
D32586 N32586 0 diode
R32587 N32586 N32587 10
D32587 N32587 0 diode
R32588 N32587 N32588 10
D32588 N32588 0 diode
R32589 N32588 N32589 10
D32589 N32589 0 diode
R32590 N32589 N32590 10
D32590 N32590 0 diode
R32591 N32590 N32591 10
D32591 N32591 0 diode
R32592 N32591 N32592 10
D32592 N32592 0 diode
R32593 N32592 N32593 10
D32593 N32593 0 diode
R32594 N32593 N32594 10
D32594 N32594 0 diode
R32595 N32594 N32595 10
D32595 N32595 0 diode
R32596 N32595 N32596 10
D32596 N32596 0 diode
R32597 N32596 N32597 10
D32597 N32597 0 diode
R32598 N32597 N32598 10
D32598 N32598 0 diode
R32599 N32598 N32599 10
D32599 N32599 0 diode
R32600 N32599 N32600 10
D32600 N32600 0 diode
R32601 N32600 N32601 10
D32601 N32601 0 diode
R32602 N32601 N32602 10
D32602 N32602 0 diode
R32603 N32602 N32603 10
D32603 N32603 0 diode
R32604 N32603 N32604 10
D32604 N32604 0 diode
R32605 N32604 N32605 10
D32605 N32605 0 diode
R32606 N32605 N32606 10
D32606 N32606 0 diode
R32607 N32606 N32607 10
D32607 N32607 0 diode
R32608 N32607 N32608 10
D32608 N32608 0 diode
R32609 N32608 N32609 10
D32609 N32609 0 diode
R32610 N32609 N32610 10
D32610 N32610 0 diode
R32611 N32610 N32611 10
D32611 N32611 0 diode
R32612 N32611 N32612 10
D32612 N32612 0 diode
R32613 N32612 N32613 10
D32613 N32613 0 diode
R32614 N32613 N32614 10
D32614 N32614 0 diode
R32615 N32614 N32615 10
D32615 N32615 0 diode
R32616 N32615 N32616 10
D32616 N32616 0 diode
R32617 N32616 N32617 10
D32617 N32617 0 diode
R32618 N32617 N32618 10
D32618 N32618 0 diode
R32619 N32618 N32619 10
D32619 N32619 0 diode
R32620 N32619 N32620 10
D32620 N32620 0 diode
R32621 N32620 N32621 10
D32621 N32621 0 diode
R32622 N32621 N32622 10
D32622 N32622 0 diode
R32623 N32622 N32623 10
D32623 N32623 0 diode
R32624 N32623 N32624 10
D32624 N32624 0 diode
R32625 N32624 N32625 10
D32625 N32625 0 diode
R32626 N32625 N32626 10
D32626 N32626 0 diode
R32627 N32626 N32627 10
D32627 N32627 0 diode
R32628 N32627 N32628 10
D32628 N32628 0 diode
R32629 N32628 N32629 10
D32629 N32629 0 diode
R32630 N32629 N32630 10
D32630 N32630 0 diode
R32631 N32630 N32631 10
D32631 N32631 0 diode
R32632 N32631 N32632 10
D32632 N32632 0 diode
R32633 N32632 N32633 10
D32633 N32633 0 diode
R32634 N32633 N32634 10
D32634 N32634 0 diode
R32635 N32634 N32635 10
D32635 N32635 0 diode
R32636 N32635 N32636 10
D32636 N32636 0 diode
R32637 N32636 N32637 10
D32637 N32637 0 diode
R32638 N32637 N32638 10
D32638 N32638 0 diode
R32639 N32638 N32639 10
D32639 N32639 0 diode
R32640 N32639 N32640 10
D32640 N32640 0 diode
R32641 N32640 N32641 10
D32641 N32641 0 diode
R32642 N32641 N32642 10
D32642 N32642 0 diode
R32643 N32642 N32643 10
D32643 N32643 0 diode
R32644 N32643 N32644 10
D32644 N32644 0 diode
R32645 N32644 N32645 10
D32645 N32645 0 diode
R32646 N32645 N32646 10
D32646 N32646 0 diode
R32647 N32646 N32647 10
D32647 N32647 0 diode
R32648 N32647 N32648 10
D32648 N32648 0 diode
R32649 N32648 N32649 10
D32649 N32649 0 diode
R32650 N32649 N32650 10
D32650 N32650 0 diode
R32651 N32650 N32651 10
D32651 N32651 0 diode
R32652 N32651 N32652 10
D32652 N32652 0 diode
R32653 N32652 N32653 10
D32653 N32653 0 diode
R32654 N32653 N32654 10
D32654 N32654 0 diode
R32655 N32654 N32655 10
D32655 N32655 0 diode
R32656 N32655 N32656 10
D32656 N32656 0 diode
R32657 N32656 N32657 10
D32657 N32657 0 diode
R32658 N32657 N32658 10
D32658 N32658 0 diode
R32659 N32658 N32659 10
D32659 N32659 0 diode
R32660 N32659 N32660 10
D32660 N32660 0 diode
R32661 N32660 N32661 10
D32661 N32661 0 diode
R32662 N32661 N32662 10
D32662 N32662 0 diode
R32663 N32662 N32663 10
D32663 N32663 0 diode
R32664 N32663 N32664 10
D32664 N32664 0 diode
R32665 N32664 N32665 10
D32665 N32665 0 diode
R32666 N32665 N32666 10
D32666 N32666 0 diode
R32667 N32666 N32667 10
D32667 N32667 0 diode
R32668 N32667 N32668 10
D32668 N32668 0 diode
R32669 N32668 N32669 10
D32669 N32669 0 diode
R32670 N32669 N32670 10
D32670 N32670 0 diode
R32671 N32670 N32671 10
D32671 N32671 0 diode
R32672 N32671 N32672 10
D32672 N32672 0 diode
R32673 N32672 N32673 10
D32673 N32673 0 diode
R32674 N32673 N32674 10
D32674 N32674 0 diode
R32675 N32674 N32675 10
D32675 N32675 0 diode
R32676 N32675 N32676 10
D32676 N32676 0 diode
R32677 N32676 N32677 10
D32677 N32677 0 diode
R32678 N32677 N32678 10
D32678 N32678 0 diode
R32679 N32678 N32679 10
D32679 N32679 0 diode
R32680 N32679 N32680 10
D32680 N32680 0 diode
R32681 N32680 N32681 10
D32681 N32681 0 diode
R32682 N32681 N32682 10
D32682 N32682 0 diode
R32683 N32682 N32683 10
D32683 N32683 0 diode
R32684 N32683 N32684 10
D32684 N32684 0 diode
R32685 N32684 N32685 10
D32685 N32685 0 diode
R32686 N32685 N32686 10
D32686 N32686 0 diode
R32687 N32686 N32687 10
D32687 N32687 0 diode
R32688 N32687 N32688 10
D32688 N32688 0 diode
R32689 N32688 N32689 10
D32689 N32689 0 diode
R32690 N32689 N32690 10
D32690 N32690 0 diode
R32691 N32690 N32691 10
D32691 N32691 0 diode
R32692 N32691 N32692 10
D32692 N32692 0 diode
R32693 N32692 N32693 10
D32693 N32693 0 diode
R32694 N32693 N32694 10
D32694 N32694 0 diode
R32695 N32694 N32695 10
D32695 N32695 0 diode
R32696 N32695 N32696 10
D32696 N32696 0 diode
R32697 N32696 N32697 10
D32697 N32697 0 diode
R32698 N32697 N32698 10
D32698 N32698 0 diode
R32699 N32698 N32699 10
D32699 N32699 0 diode
R32700 N32699 N32700 10
D32700 N32700 0 diode
R32701 N32700 N32701 10
D32701 N32701 0 diode
R32702 N32701 N32702 10
D32702 N32702 0 diode
R32703 N32702 N32703 10
D32703 N32703 0 diode
R32704 N32703 N32704 10
D32704 N32704 0 diode
R32705 N32704 N32705 10
D32705 N32705 0 diode
R32706 N32705 N32706 10
D32706 N32706 0 diode
R32707 N32706 N32707 10
D32707 N32707 0 diode
R32708 N32707 N32708 10
D32708 N32708 0 diode
R32709 N32708 N32709 10
D32709 N32709 0 diode
R32710 N32709 N32710 10
D32710 N32710 0 diode
R32711 N32710 N32711 10
D32711 N32711 0 diode
R32712 N32711 N32712 10
D32712 N32712 0 diode
R32713 N32712 N32713 10
D32713 N32713 0 diode
R32714 N32713 N32714 10
D32714 N32714 0 diode
R32715 N32714 N32715 10
D32715 N32715 0 diode
R32716 N32715 N32716 10
D32716 N32716 0 diode
R32717 N32716 N32717 10
D32717 N32717 0 diode
R32718 N32717 N32718 10
D32718 N32718 0 diode
R32719 N32718 N32719 10
D32719 N32719 0 diode
R32720 N32719 N32720 10
D32720 N32720 0 diode
R32721 N32720 N32721 10
D32721 N32721 0 diode
R32722 N32721 N32722 10
D32722 N32722 0 diode
R32723 N32722 N32723 10
D32723 N32723 0 diode
R32724 N32723 N32724 10
D32724 N32724 0 diode
R32725 N32724 N32725 10
D32725 N32725 0 diode
R32726 N32725 N32726 10
D32726 N32726 0 diode
R32727 N32726 N32727 10
D32727 N32727 0 diode
R32728 N32727 N32728 10
D32728 N32728 0 diode
R32729 N32728 N32729 10
D32729 N32729 0 diode
R32730 N32729 N32730 10
D32730 N32730 0 diode
R32731 N32730 N32731 10
D32731 N32731 0 diode
R32732 N32731 N32732 10
D32732 N32732 0 diode
R32733 N32732 N32733 10
D32733 N32733 0 diode
R32734 N32733 N32734 10
D32734 N32734 0 diode
R32735 N32734 N32735 10
D32735 N32735 0 diode
R32736 N32735 N32736 10
D32736 N32736 0 diode
R32737 N32736 N32737 10
D32737 N32737 0 diode
R32738 N32737 N32738 10
D32738 N32738 0 diode
R32739 N32738 N32739 10
D32739 N32739 0 diode
R32740 N32739 N32740 10
D32740 N32740 0 diode
R32741 N32740 N32741 10
D32741 N32741 0 diode
R32742 N32741 N32742 10
D32742 N32742 0 diode
R32743 N32742 N32743 10
D32743 N32743 0 diode
R32744 N32743 N32744 10
D32744 N32744 0 diode
R32745 N32744 N32745 10
D32745 N32745 0 diode
R32746 N32745 N32746 10
D32746 N32746 0 diode
R32747 N32746 N32747 10
D32747 N32747 0 diode
R32748 N32747 N32748 10
D32748 N32748 0 diode
R32749 N32748 N32749 10
D32749 N32749 0 diode
R32750 N32749 N32750 10
D32750 N32750 0 diode
R32751 N32750 N32751 10
D32751 N32751 0 diode
R32752 N32751 N32752 10
D32752 N32752 0 diode
R32753 N32752 N32753 10
D32753 N32753 0 diode
R32754 N32753 N32754 10
D32754 N32754 0 diode
R32755 N32754 N32755 10
D32755 N32755 0 diode
R32756 N32755 N32756 10
D32756 N32756 0 diode
R32757 N32756 N32757 10
D32757 N32757 0 diode
R32758 N32757 N32758 10
D32758 N32758 0 diode
R32759 N32758 N32759 10
D32759 N32759 0 diode
R32760 N32759 N32760 10
D32760 N32760 0 diode
R32761 N32760 N32761 10
D32761 N32761 0 diode
R32762 N32761 N32762 10
D32762 N32762 0 diode
R32763 N32762 N32763 10
D32763 N32763 0 diode
R32764 N32763 N32764 10
D32764 N32764 0 diode
R32765 N32764 N32765 10
D32765 N32765 0 diode
R32766 N32765 N32766 10
D32766 N32766 0 diode
R32767 N32766 N32767 10
D32767 N32767 0 diode
R32768 N32767 N32768 10
D32768 N32768 0 diode
R32769 N32768 N32769 10
D32769 N32769 0 diode
R32770 N32769 N32770 10
D32770 N32770 0 diode
R32771 N32770 N32771 10
D32771 N32771 0 diode
R32772 N32771 N32772 10
D32772 N32772 0 diode
R32773 N32772 N32773 10
D32773 N32773 0 diode
R32774 N32773 N32774 10
D32774 N32774 0 diode
R32775 N32774 N32775 10
D32775 N32775 0 diode
R32776 N32775 N32776 10
D32776 N32776 0 diode
R32777 N32776 N32777 10
D32777 N32777 0 diode
R32778 N32777 N32778 10
D32778 N32778 0 diode
R32779 N32778 N32779 10
D32779 N32779 0 diode
R32780 N32779 N32780 10
D32780 N32780 0 diode
R32781 N32780 N32781 10
D32781 N32781 0 diode
R32782 N32781 N32782 10
D32782 N32782 0 diode
R32783 N32782 N32783 10
D32783 N32783 0 diode
R32784 N32783 N32784 10
D32784 N32784 0 diode
R32785 N32784 N32785 10
D32785 N32785 0 diode
R32786 N32785 N32786 10
D32786 N32786 0 diode
R32787 N32786 N32787 10
D32787 N32787 0 diode
R32788 N32787 N32788 10
D32788 N32788 0 diode
R32789 N32788 N32789 10
D32789 N32789 0 diode
R32790 N32789 N32790 10
D32790 N32790 0 diode
R32791 N32790 N32791 10
D32791 N32791 0 diode
R32792 N32791 N32792 10
D32792 N32792 0 diode
R32793 N32792 N32793 10
D32793 N32793 0 diode
R32794 N32793 N32794 10
D32794 N32794 0 diode
R32795 N32794 N32795 10
D32795 N32795 0 diode
R32796 N32795 N32796 10
D32796 N32796 0 diode
R32797 N32796 N32797 10
D32797 N32797 0 diode
R32798 N32797 N32798 10
D32798 N32798 0 diode
R32799 N32798 N32799 10
D32799 N32799 0 diode
R32800 N32799 N32800 10
D32800 N32800 0 diode
R32801 N32800 N32801 10
D32801 N32801 0 diode
R32802 N32801 N32802 10
D32802 N32802 0 diode
R32803 N32802 N32803 10
D32803 N32803 0 diode
R32804 N32803 N32804 10
D32804 N32804 0 diode
R32805 N32804 N32805 10
D32805 N32805 0 diode
R32806 N32805 N32806 10
D32806 N32806 0 diode
R32807 N32806 N32807 10
D32807 N32807 0 diode
R32808 N32807 N32808 10
D32808 N32808 0 diode
R32809 N32808 N32809 10
D32809 N32809 0 diode
R32810 N32809 N32810 10
D32810 N32810 0 diode
R32811 N32810 N32811 10
D32811 N32811 0 diode
R32812 N32811 N32812 10
D32812 N32812 0 diode
R32813 N32812 N32813 10
D32813 N32813 0 diode
R32814 N32813 N32814 10
D32814 N32814 0 diode
R32815 N32814 N32815 10
D32815 N32815 0 diode
R32816 N32815 N32816 10
D32816 N32816 0 diode
R32817 N32816 N32817 10
D32817 N32817 0 diode
R32818 N32817 N32818 10
D32818 N32818 0 diode
R32819 N32818 N32819 10
D32819 N32819 0 diode
R32820 N32819 N32820 10
D32820 N32820 0 diode
R32821 N32820 N32821 10
D32821 N32821 0 diode
R32822 N32821 N32822 10
D32822 N32822 0 diode
R32823 N32822 N32823 10
D32823 N32823 0 diode
R32824 N32823 N32824 10
D32824 N32824 0 diode
R32825 N32824 N32825 10
D32825 N32825 0 diode
R32826 N32825 N32826 10
D32826 N32826 0 diode
R32827 N32826 N32827 10
D32827 N32827 0 diode
R32828 N32827 N32828 10
D32828 N32828 0 diode
R32829 N32828 N32829 10
D32829 N32829 0 diode
R32830 N32829 N32830 10
D32830 N32830 0 diode
R32831 N32830 N32831 10
D32831 N32831 0 diode
R32832 N32831 N32832 10
D32832 N32832 0 diode
R32833 N32832 N32833 10
D32833 N32833 0 diode
R32834 N32833 N32834 10
D32834 N32834 0 diode
R32835 N32834 N32835 10
D32835 N32835 0 diode
R32836 N32835 N32836 10
D32836 N32836 0 diode
R32837 N32836 N32837 10
D32837 N32837 0 diode
R32838 N32837 N32838 10
D32838 N32838 0 diode
R32839 N32838 N32839 10
D32839 N32839 0 diode
R32840 N32839 N32840 10
D32840 N32840 0 diode
R32841 N32840 N32841 10
D32841 N32841 0 diode
R32842 N32841 N32842 10
D32842 N32842 0 diode
R32843 N32842 N32843 10
D32843 N32843 0 diode
R32844 N32843 N32844 10
D32844 N32844 0 diode
R32845 N32844 N32845 10
D32845 N32845 0 diode
R32846 N32845 N32846 10
D32846 N32846 0 diode
R32847 N32846 N32847 10
D32847 N32847 0 diode
R32848 N32847 N32848 10
D32848 N32848 0 diode
R32849 N32848 N32849 10
D32849 N32849 0 diode
R32850 N32849 N32850 10
D32850 N32850 0 diode
R32851 N32850 N32851 10
D32851 N32851 0 diode
R32852 N32851 N32852 10
D32852 N32852 0 diode
R32853 N32852 N32853 10
D32853 N32853 0 diode
R32854 N32853 N32854 10
D32854 N32854 0 diode
R32855 N32854 N32855 10
D32855 N32855 0 diode
R32856 N32855 N32856 10
D32856 N32856 0 diode
R32857 N32856 N32857 10
D32857 N32857 0 diode
R32858 N32857 N32858 10
D32858 N32858 0 diode
R32859 N32858 N32859 10
D32859 N32859 0 diode
R32860 N32859 N32860 10
D32860 N32860 0 diode
R32861 N32860 N32861 10
D32861 N32861 0 diode
R32862 N32861 N32862 10
D32862 N32862 0 diode
R32863 N32862 N32863 10
D32863 N32863 0 diode
R32864 N32863 N32864 10
D32864 N32864 0 diode
R32865 N32864 N32865 10
D32865 N32865 0 diode
R32866 N32865 N32866 10
D32866 N32866 0 diode
R32867 N32866 N32867 10
D32867 N32867 0 diode
R32868 N32867 N32868 10
D32868 N32868 0 diode
R32869 N32868 N32869 10
D32869 N32869 0 diode
R32870 N32869 N32870 10
D32870 N32870 0 diode
R32871 N32870 N32871 10
D32871 N32871 0 diode
R32872 N32871 N32872 10
D32872 N32872 0 diode
R32873 N32872 N32873 10
D32873 N32873 0 diode
R32874 N32873 N32874 10
D32874 N32874 0 diode
R32875 N32874 N32875 10
D32875 N32875 0 diode
R32876 N32875 N32876 10
D32876 N32876 0 diode
R32877 N32876 N32877 10
D32877 N32877 0 diode
R32878 N32877 N32878 10
D32878 N32878 0 diode
R32879 N32878 N32879 10
D32879 N32879 0 diode
R32880 N32879 N32880 10
D32880 N32880 0 diode
R32881 N32880 N32881 10
D32881 N32881 0 diode
R32882 N32881 N32882 10
D32882 N32882 0 diode
R32883 N32882 N32883 10
D32883 N32883 0 diode
R32884 N32883 N32884 10
D32884 N32884 0 diode
R32885 N32884 N32885 10
D32885 N32885 0 diode
R32886 N32885 N32886 10
D32886 N32886 0 diode
R32887 N32886 N32887 10
D32887 N32887 0 diode
R32888 N32887 N32888 10
D32888 N32888 0 diode
R32889 N32888 N32889 10
D32889 N32889 0 diode
R32890 N32889 N32890 10
D32890 N32890 0 diode
R32891 N32890 N32891 10
D32891 N32891 0 diode
R32892 N32891 N32892 10
D32892 N32892 0 diode
R32893 N32892 N32893 10
D32893 N32893 0 diode
R32894 N32893 N32894 10
D32894 N32894 0 diode
R32895 N32894 N32895 10
D32895 N32895 0 diode
R32896 N32895 N32896 10
D32896 N32896 0 diode
R32897 N32896 N32897 10
D32897 N32897 0 diode
R32898 N32897 N32898 10
D32898 N32898 0 diode
R32899 N32898 N32899 10
D32899 N32899 0 diode
R32900 N32899 N32900 10
D32900 N32900 0 diode
R32901 N32900 N32901 10
D32901 N32901 0 diode
R32902 N32901 N32902 10
D32902 N32902 0 diode
R32903 N32902 N32903 10
D32903 N32903 0 diode
R32904 N32903 N32904 10
D32904 N32904 0 diode
R32905 N32904 N32905 10
D32905 N32905 0 diode
R32906 N32905 N32906 10
D32906 N32906 0 diode
R32907 N32906 N32907 10
D32907 N32907 0 diode
R32908 N32907 N32908 10
D32908 N32908 0 diode
R32909 N32908 N32909 10
D32909 N32909 0 diode
R32910 N32909 N32910 10
D32910 N32910 0 diode
R32911 N32910 N32911 10
D32911 N32911 0 diode
R32912 N32911 N32912 10
D32912 N32912 0 diode
R32913 N32912 N32913 10
D32913 N32913 0 diode
R32914 N32913 N32914 10
D32914 N32914 0 diode
R32915 N32914 N32915 10
D32915 N32915 0 diode
R32916 N32915 N32916 10
D32916 N32916 0 diode
R32917 N32916 N32917 10
D32917 N32917 0 diode
R32918 N32917 N32918 10
D32918 N32918 0 diode
R32919 N32918 N32919 10
D32919 N32919 0 diode
R32920 N32919 N32920 10
D32920 N32920 0 diode
R32921 N32920 N32921 10
D32921 N32921 0 diode
R32922 N32921 N32922 10
D32922 N32922 0 diode
R32923 N32922 N32923 10
D32923 N32923 0 diode
R32924 N32923 N32924 10
D32924 N32924 0 diode
R32925 N32924 N32925 10
D32925 N32925 0 diode
R32926 N32925 N32926 10
D32926 N32926 0 diode
R32927 N32926 N32927 10
D32927 N32927 0 diode
R32928 N32927 N32928 10
D32928 N32928 0 diode
R32929 N32928 N32929 10
D32929 N32929 0 diode
R32930 N32929 N32930 10
D32930 N32930 0 diode
R32931 N32930 N32931 10
D32931 N32931 0 diode
R32932 N32931 N32932 10
D32932 N32932 0 diode
R32933 N32932 N32933 10
D32933 N32933 0 diode
R32934 N32933 N32934 10
D32934 N32934 0 diode
R32935 N32934 N32935 10
D32935 N32935 0 diode
R32936 N32935 N32936 10
D32936 N32936 0 diode
R32937 N32936 N32937 10
D32937 N32937 0 diode
R32938 N32937 N32938 10
D32938 N32938 0 diode
R32939 N32938 N32939 10
D32939 N32939 0 diode
R32940 N32939 N32940 10
D32940 N32940 0 diode
R32941 N32940 N32941 10
D32941 N32941 0 diode
R32942 N32941 N32942 10
D32942 N32942 0 diode
R32943 N32942 N32943 10
D32943 N32943 0 diode
R32944 N32943 N32944 10
D32944 N32944 0 diode
R32945 N32944 N32945 10
D32945 N32945 0 diode
R32946 N32945 N32946 10
D32946 N32946 0 diode
R32947 N32946 N32947 10
D32947 N32947 0 diode
R32948 N32947 N32948 10
D32948 N32948 0 diode
R32949 N32948 N32949 10
D32949 N32949 0 diode
R32950 N32949 N32950 10
D32950 N32950 0 diode
R32951 N32950 N32951 10
D32951 N32951 0 diode
R32952 N32951 N32952 10
D32952 N32952 0 diode
R32953 N32952 N32953 10
D32953 N32953 0 diode
R32954 N32953 N32954 10
D32954 N32954 0 diode
R32955 N32954 N32955 10
D32955 N32955 0 diode
R32956 N32955 N32956 10
D32956 N32956 0 diode
R32957 N32956 N32957 10
D32957 N32957 0 diode
R32958 N32957 N32958 10
D32958 N32958 0 diode
R32959 N32958 N32959 10
D32959 N32959 0 diode
R32960 N32959 N32960 10
D32960 N32960 0 diode
R32961 N32960 N32961 10
D32961 N32961 0 diode
R32962 N32961 N32962 10
D32962 N32962 0 diode
R32963 N32962 N32963 10
D32963 N32963 0 diode
R32964 N32963 N32964 10
D32964 N32964 0 diode
R32965 N32964 N32965 10
D32965 N32965 0 diode
R32966 N32965 N32966 10
D32966 N32966 0 diode
R32967 N32966 N32967 10
D32967 N32967 0 diode
R32968 N32967 N32968 10
D32968 N32968 0 diode
R32969 N32968 N32969 10
D32969 N32969 0 diode
R32970 N32969 N32970 10
D32970 N32970 0 diode
R32971 N32970 N32971 10
D32971 N32971 0 diode
R32972 N32971 N32972 10
D32972 N32972 0 diode
R32973 N32972 N32973 10
D32973 N32973 0 diode
R32974 N32973 N32974 10
D32974 N32974 0 diode
R32975 N32974 N32975 10
D32975 N32975 0 diode
R32976 N32975 N32976 10
D32976 N32976 0 diode
R32977 N32976 N32977 10
D32977 N32977 0 diode
R32978 N32977 N32978 10
D32978 N32978 0 diode
R32979 N32978 N32979 10
D32979 N32979 0 diode
R32980 N32979 N32980 10
D32980 N32980 0 diode
R32981 N32980 N32981 10
D32981 N32981 0 diode
R32982 N32981 N32982 10
D32982 N32982 0 diode
R32983 N32982 N32983 10
D32983 N32983 0 diode
R32984 N32983 N32984 10
D32984 N32984 0 diode
R32985 N32984 N32985 10
D32985 N32985 0 diode
R32986 N32985 N32986 10
D32986 N32986 0 diode
R32987 N32986 N32987 10
D32987 N32987 0 diode
R32988 N32987 N32988 10
D32988 N32988 0 diode
R32989 N32988 N32989 10
D32989 N32989 0 diode
R32990 N32989 N32990 10
D32990 N32990 0 diode
R32991 N32990 N32991 10
D32991 N32991 0 diode
R32992 N32991 N32992 10
D32992 N32992 0 diode
R32993 N32992 N32993 10
D32993 N32993 0 diode
R32994 N32993 N32994 10
D32994 N32994 0 diode
R32995 N32994 N32995 10
D32995 N32995 0 diode
R32996 N32995 N32996 10
D32996 N32996 0 diode
R32997 N32996 N32997 10
D32997 N32997 0 diode
R32998 N32997 N32998 10
D32998 N32998 0 diode
R32999 N32998 N32999 10
D32999 N32999 0 diode
R33000 N32999 N33000 10
D33000 N33000 0 diode
R33001 N33000 N33001 10
D33001 N33001 0 diode
R33002 N33001 N33002 10
D33002 N33002 0 diode
R33003 N33002 N33003 10
D33003 N33003 0 diode
R33004 N33003 N33004 10
D33004 N33004 0 diode
R33005 N33004 N33005 10
D33005 N33005 0 diode
R33006 N33005 N33006 10
D33006 N33006 0 diode
R33007 N33006 N33007 10
D33007 N33007 0 diode
R33008 N33007 N33008 10
D33008 N33008 0 diode
R33009 N33008 N33009 10
D33009 N33009 0 diode
R33010 N33009 N33010 10
D33010 N33010 0 diode
R33011 N33010 N33011 10
D33011 N33011 0 diode
R33012 N33011 N33012 10
D33012 N33012 0 diode
R33013 N33012 N33013 10
D33013 N33013 0 diode
R33014 N33013 N33014 10
D33014 N33014 0 diode
R33015 N33014 N33015 10
D33015 N33015 0 diode
R33016 N33015 N33016 10
D33016 N33016 0 diode
R33017 N33016 N33017 10
D33017 N33017 0 diode
R33018 N33017 N33018 10
D33018 N33018 0 diode
R33019 N33018 N33019 10
D33019 N33019 0 diode
R33020 N33019 N33020 10
D33020 N33020 0 diode
R33021 N33020 N33021 10
D33021 N33021 0 diode
R33022 N33021 N33022 10
D33022 N33022 0 diode
R33023 N33022 N33023 10
D33023 N33023 0 diode
R33024 N33023 N33024 10
D33024 N33024 0 diode
R33025 N33024 N33025 10
D33025 N33025 0 diode
R33026 N33025 N33026 10
D33026 N33026 0 diode
R33027 N33026 N33027 10
D33027 N33027 0 diode
R33028 N33027 N33028 10
D33028 N33028 0 diode
R33029 N33028 N33029 10
D33029 N33029 0 diode
R33030 N33029 N33030 10
D33030 N33030 0 diode
R33031 N33030 N33031 10
D33031 N33031 0 diode
R33032 N33031 N33032 10
D33032 N33032 0 diode
R33033 N33032 N33033 10
D33033 N33033 0 diode
R33034 N33033 N33034 10
D33034 N33034 0 diode
R33035 N33034 N33035 10
D33035 N33035 0 diode
R33036 N33035 N33036 10
D33036 N33036 0 diode
R33037 N33036 N33037 10
D33037 N33037 0 diode
R33038 N33037 N33038 10
D33038 N33038 0 diode
R33039 N33038 N33039 10
D33039 N33039 0 diode
R33040 N33039 N33040 10
D33040 N33040 0 diode
R33041 N33040 N33041 10
D33041 N33041 0 diode
R33042 N33041 N33042 10
D33042 N33042 0 diode
R33043 N33042 N33043 10
D33043 N33043 0 diode
R33044 N33043 N33044 10
D33044 N33044 0 diode
R33045 N33044 N33045 10
D33045 N33045 0 diode
R33046 N33045 N33046 10
D33046 N33046 0 diode
R33047 N33046 N33047 10
D33047 N33047 0 diode
R33048 N33047 N33048 10
D33048 N33048 0 diode
R33049 N33048 N33049 10
D33049 N33049 0 diode
R33050 N33049 N33050 10
D33050 N33050 0 diode
R33051 N33050 N33051 10
D33051 N33051 0 diode
R33052 N33051 N33052 10
D33052 N33052 0 diode
R33053 N33052 N33053 10
D33053 N33053 0 diode
R33054 N33053 N33054 10
D33054 N33054 0 diode
R33055 N33054 N33055 10
D33055 N33055 0 diode
R33056 N33055 N33056 10
D33056 N33056 0 diode
R33057 N33056 N33057 10
D33057 N33057 0 diode
R33058 N33057 N33058 10
D33058 N33058 0 diode
R33059 N33058 N33059 10
D33059 N33059 0 diode
R33060 N33059 N33060 10
D33060 N33060 0 diode
R33061 N33060 N33061 10
D33061 N33061 0 diode
R33062 N33061 N33062 10
D33062 N33062 0 diode
R33063 N33062 N33063 10
D33063 N33063 0 diode
R33064 N33063 N33064 10
D33064 N33064 0 diode
R33065 N33064 N33065 10
D33065 N33065 0 diode
R33066 N33065 N33066 10
D33066 N33066 0 diode
R33067 N33066 N33067 10
D33067 N33067 0 diode
R33068 N33067 N33068 10
D33068 N33068 0 diode
R33069 N33068 N33069 10
D33069 N33069 0 diode
R33070 N33069 N33070 10
D33070 N33070 0 diode
R33071 N33070 N33071 10
D33071 N33071 0 diode
R33072 N33071 N33072 10
D33072 N33072 0 diode
R33073 N33072 N33073 10
D33073 N33073 0 diode
R33074 N33073 N33074 10
D33074 N33074 0 diode
R33075 N33074 N33075 10
D33075 N33075 0 diode
R33076 N33075 N33076 10
D33076 N33076 0 diode
R33077 N33076 N33077 10
D33077 N33077 0 diode
R33078 N33077 N33078 10
D33078 N33078 0 diode
R33079 N33078 N33079 10
D33079 N33079 0 diode
R33080 N33079 N33080 10
D33080 N33080 0 diode
R33081 N33080 N33081 10
D33081 N33081 0 diode
R33082 N33081 N33082 10
D33082 N33082 0 diode
R33083 N33082 N33083 10
D33083 N33083 0 diode
R33084 N33083 N33084 10
D33084 N33084 0 diode
R33085 N33084 N33085 10
D33085 N33085 0 diode
R33086 N33085 N33086 10
D33086 N33086 0 diode
R33087 N33086 N33087 10
D33087 N33087 0 diode
R33088 N33087 N33088 10
D33088 N33088 0 diode
R33089 N33088 N33089 10
D33089 N33089 0 diode
R33090 N33089 N33090 10
D33090 N33090 0 diode
R33091 N33090 N33091 10
D33091 N33091 0 diode
R33092 N33091 N33092 10
D33092 N33092 0 diode
R33093 N33092 N33093 10
D33093 N33093 0 diode
R33094 N33093 N33094 10
D33094 N33094 0 diode
R33095 N33094 N33095 10
D33095 N33095 0 diode
R33096 N33095 N33096 10
D33096 N33096 0 diode
R33097 N33096 N33097 10
D33097 N33097 0 diode
R33098 N33097 N33098 10
D33098 N33098 0 diode
R33099 N33098 N33099 10
D33099 N33099 0 diode
R33100 N33099 N33100 10
D33100 N33100 0 diode
R33101 N33100 N33101 10
D33101 N33101 0 diode
R33102 N33101 N33102 10
D33102 N33102 0 diode
R33103 N33102 N33103 10
D33103 N33103 0 diode
R33104 N33103 N33104 10
D33104 N33104 0 diode
R33105 N33104 N33105 10
D33105 N33105 0 diode
R33106 N33105 N33106 10
D33106 N33106 0 diode
R33107 N33106 N33107 10
D33107 N33107 0 diode
R33108 N33107 N33108 10
D33108 N33108 0 diode
R33109 N33108 N33109 10
D33109 N33109 0 diode
R33110 N33109 N33110 10
D33110 N33110 0 diode
R33111 N33110 N33111 10
D33111 N33111 0 diode
R33112 N33111 N33112 10
D33112 N33112 0 diode
R33113 N33112 N33113 10
D33113 N33113 0 diode
R33114 N33113 N33114 10
D33114 N33114 0 diode
R33115 N33114 N33115 10
D33115 N33115 0 diode
R33116 N33115 N33116 10
D33116 N33116 0 diode
R33117 N33116 N33117 10
D33117 N33117 0 diode
R33118 N33117 N33118 10
D33118 N33118 0 diode
R33119 N33118 N33119 10
D33119 N33119 0 diode
R33120 N33119 N33120 10
D33120 N33120 0 diode
R33121 N33120 N33121 10
D33121 N33121 0 diode
R33122 N33121 N33122 10
D33122 N33122 0 diode
R33123 N33122 N33123 10
D33123 N33123 0 diode
R33124 N33123 N33124 10
D33124 N33124 0 diode
R33125 N33124 N33125 10
D33125 N33125 0 diode
R33126 N33125 N33126 10
D33126 N33126 0 diode
R33127 N33126 N33127 10
D33127 N33127 0 diode
R33128 N33127 N33128 10
D33128 N33128 0 diode
R33129 N33128 N33129 10
D33129 N33129 0 diode
R33130 N33129 N33130 10
D33130 N33130 0 diode
R33131 N33130 N33131 10
D33131 N33131 0 diode
R33132 N33131 N33132 10
D33132 N33132 0 diode
R33133 N33132 N33133 10
D33133 N33133 0 diode
R33134 N33133 N33134 10
D33134 N33134 0 diode
R33135 N33134 N33135 10
D33135 N33135 0 diode
R33136 N33135 N33136 10
D33136 N33136 0 diode
R33137 N33136 N33137 10
D33137 N33137 0 diode
R33138 N33137 N33138 10
D33138 N33138 0 diode
R33139 N33138 N33139 10
D33139 N33139 0 diode
R33140 N33139 N33140 10
D33140 N33140 0 diode
R33141 N33140 N33141 10
D33141 N33141 0 diode
R33142 N33141 N33142 10
D33142 N33142 0 diode
R33143 N33142 N33143 10
D33143 N33143 0 diode
R33144 N33143 N33144 10
D33144 N33144 0 diode
R33145 N33144 N33145 10
D33145 N33145 0 diode
R33146 N33145 N33146 10
D33146 N33146 0 diode
R33147 N33146 N33147 10
D33147 N33147 0 diode
R33148 N33147 N33148 10
D33148 N33148 0 diode
R33149 N33148 N33149 10
D33149 N33149 0 diode
R33150 N33149 N33150 10
D33150 N33150 0 diode
R33151 N33150 N33151 10
D33151 N33151 0 diode
R33152 N33151 N33152 10
D33152 N33152 0 diode
R33153 N33152 N33153 10
D33153 N33153 0 diode
R33154 N33153 N33154 10
D33154 N33154 0 diode
R33155 N33154 N33155 10
D33155 N33155 0 diode
R33156 N33155 N33156 10
D33156 N33156 0 diode
R33157 N33156 N33157 10
D33157 N33157 0 diode
R33158 N33157 N33158 10
D33158 N33158 0 diode
R33159 N33158 N33159 10
D33159 N33159 0 diode
R33160 N33159 N33160 10
D33160 N33160 0 diode
R33161 N33160 N33161 10
D33161 N33161 0 diode
R33162 N33161 N33162 10
D33162 N33162 0 diode
R33163 N33162 N33163 10
D33163 N33163 0 diode
R33164 N33163 N33164 10
D33164 N33164 0 diode
R33165 N33164 N33165 10
D33165 N33165 0 diode
R33166 N33165 N33166 10
D33166 N33166 0 diode
R33167 N33166 N33167 10
D33167 N33167 0 diode
R33168 N33167 N33168 10
D33168 N33168 0 diode
R33169 N33168 N33169 10
D33169 N33169 0 diode
R33170 N33169 N33170 10
D33170 N33170 0 diode
R33171 N33170 N33171 10
D33171 N33171 0 diode
R33172 N33171 N33172 10
D33172 N33172 0 diode
R33173 N33172 N33173 10
D33173 N33173 0 diode
R33174 N33173 N33174 10
D33174 N33174 0 diode
R33175 N33174 N33175 10
D33175 N33175 0 diode
R33176 N33175 N33176 10
D33176 N33176 0 diode
R33177 N33176 N33177 10
D33177 N33177 0 diode
R33178 N33177 N33178 10
D33178 N33178 0 diode
R33179 N33178 N33179 10
D33179 N33179 0 diode
R33180 N33179 N33180 10
D33180 N33180 0 diode
R33181 N33180 N33181 10
D33181 N33181 0 diode
R33182 N33181 N33182 10
D33182 N33182 0 diode
R33183 N33182 N33183 10
D33183 N33183 0 diode
R33184 N33183 N33184 10
D33184 N33184 0 diode
R33185 N33184 N33185 10
D33185 N33185 0 diode
R33186 N33185 N33186 10
D33186 N33186 0 diode
R33187 N33186 N33187 10
D33187 N33187 0 diode
R33188 N33187 N33188 10
D33188 N33188 0 diode
R33189 N33188 N33189 10
D33189 N33189 0 diode
R33190 N33189 N33190 10
D33190 N33190 0 diode
R33191 N33190 N33191 10
D33191 N33191 0 diode
R33192 N33191 N33192 10
D33192 N33192 0 diode
R33193 N33192 N33193 10
D33193 N33193 0 diode
R33194 N33193 N33194 10
D33194 N33194 0 diode
R33195 N33194 N33195 10
D33195 N33195 0 diode
R33196 N33195 N33196 10
D33196 N33196 0 diode
R33197 N33196 N33197 10
D33197 N33197 0 diode
R33198 N33197 N33198 10
D33198 N33198 0 diode
R33199 N33198 N33199 10
D33199 N33199 0 diode
R33200 N33199 N33200 10
D33200 N33200 0 diode
R33201 N33200 N33201 10
D33201 N33201 0 diode
R33202 N33201 N33202 10
D33202 N33202 0 diode
R33203 N33202 N33203 10
D33203 N33203 0 diode
R33204 N33203 N33204 10
D33204 N33204 0 diode
R33205 N33204 N33205 10
D33205 N33205 0 diode
R33206 N33205 N33206 10
D33206 N33206 0 diode
R33207 N33206 N33207 10
D33207 N33207 0 diode
R33208 N33207 N33208 10
D33208 N33208 0 diode
R33209 N33208 N33209 10
D33209 N33209 0 diode
R33210 N33209 N33210 10
D33210 N33210 0 diode
R33211 N33210 N33211 10
D33211 N33211 0 diode
R33212 N33211 N33212 10
D33212 N33212 0 diode
R33213 N33212 N33213 10
D33213 N33213 0 diode
R33214 N33213 N33214 10
D33214 N33214 0 diode
R33215 N33214 N33215 10
D33215 N33215 0 diode
R33216 N33215 N33216 10
D33216 N33216 0 diode
R33217 N33216 N33217 10
D33217 N33217 0 diode
R33218 N33217 N33218 10
D33218 N33218 0 diode
R33219 N33218 N33219 10
D33219 N33219 0 diode
R33220 N33219 N33220 10
D33220 N33220 0 diode
R33221 N33220 N33221 10
D33221 N33221 0 diode
R33222 N33221 N33222 10
D33222 N33222 0 diode
R33223 N33222 N33223 10
D33223 N33223 0 diode
R33224 N33223 N33224 10
D33224 N33224 0 diode
R33225 N33224 N33225 10
D33225 N33225 0 diode
R33226 N33225 N33226 10
D33226 N33226 0 diode
R33227 N33226 N33227 10
D33227 N33227 0 diode
R33228 N33227 N33228 10
D33228 N33228 0 diode
R33229 N33228 N33229 10
D33229 N33229 0 diode
R33230 N33229 N33230 10
D33230 N33230 0 diode
R33231 N33230 N33231 10
D33231 N33231 0 diode
R33232 N33231 N33232 10
D33232 N33232 0 diode
R33233 N33232 N33233 10
D33233 N33233 0 diode
R33234 N33233 N33234 10
D33234 N33234 0 diode
R33235 N33234 N33235 10
D33235 N33235 0 diode
R33236 N33235 N33236 10
D33236 N33236 0 diode
R33237 N33236 N33237 10
D33237 N33237 0 diode
R33238 N33237 N33238 10
D33238 N33238 0 diode
R33239 N33238 N33239 10
D33239 N33239 0 diode
R33240 N33239 N33240 10
D33240 N33240 0 diode
R33241 N33240 N33241 10
D33241 N33241 0 diode
R33242 N33241 N33242 10
D33242 N33242 0 diode
R33243 N33242 N33243 10
D33243 N33243 0 diode
R33244 N33243 N33244 10
D33244 N33244 0 diode
R33245 N33244 N33245 10
D33245 N33245 0 diode
R33246 N33245 N33246 10
D33246 N33246 0 diode
R33247 N33246 N33247 10
D33247 N33247 0 diode
R33248 N33247 N33248 10
D33248 N33248 0 diode
R33249 N33248 N33249 10
D33249 N33249 0 diode
R33250 N33249 N33250 10
D33250 N33250 0 diode
R33251 N33250 N33251 10
D33251 N33251 0 diode
R33252 N33251 N33252 10
D33252 N33252 0 diode
R33253 N33252 N33253 10
D33253 N33253 0 diode
R33254 N33253 N33254 10
D33254 N33254 0 diode
R33255 N33254 N33255 10
D33255 N33255 0 diode
R33256 N33255 N33256 10
D33256 N33256 0 diode
R33257 N33256 N33257 10
D33257 N33257 0 diode
R33258 N33257 N33258 10
D33258 N33258 0 diode
R33259 N33258 N33259 10
D33259 N33259 0 diode
R33260 N33259 N33260 10
D33260 N33260 0 diode
R33261 N33260 N33261 10
D33261 N33261 0 diode
R33262 N33261 N33262 10
D33262 N33262 0 diode
R33263 N33262 N33263 10
D33263 N33263 0 diode
R33264 N33263 N33264 10
D33264 N33264 0 diode
R33265 N33264 N33265 10
D33265 N33265 0 diode
R33266 N33265 N33266 10
D33266 N33266 0 diode
R33267 N33266 N33267 10
D33267 N33267 0 diode
R33268 N33267 N33268 10
D33268 N33268 0 diode
R33269 N33268 N33269 10
D33269 N33269 0 diode
R33270 N33269 N33270 10
D33270 N33270 0 diode
R33271 N33270 N33271 10
D33271 N33271 0 diode
R33272 N33271 N33272 10
D33272 N33272 0 diode
R33273 N33272 N33273 10
D33273 N33273 0 diode
R33274 N33273 N33274 10
D33274 N33274 0 diode
R33275 N33274 N33275 10
D33275 N33275 0 diode
R33276 N33275 N33276 10
D33276 N33276 0 diode
R33277 N33276 N33277 10
D33277 N33277 0 diode
R33278 N33277 N33278 10
D33278 N33278 0 diode
R33279 N33278 N33279 10
D33279 N33279 0 diode
R33280 N33279 N33280 10
D33280 N33280 0 diode
R33281 N33280 N33281 10
D33281 N33281 0 diode
R33282 N33281 N33282 10
D33282 N33282 0 diode
R33283 N33282 N33283 10
D33283 N33283 0 diode
R33284 N33283 N33284 10
D33284 N33284 0 diode
R33285 N33284 N33285 10
D33285 N33285 0 diode
R33286 N33285 N33286 10
D33286 N33286 0 diode
R33287 N33286 N33287 10
D33287 N33287 0 diode
R33288 N33287 N33288 10
D33288 N33288 0 diode
R33289 N33288 N33289 10
D33289 N33289 0 diode
R33290 N33289 N33290 10
D33290 N33290 0 diode
R33291 N33290 N33291 10
D33291 N33291 0 diode
R33292 N33291 N33292 10
D33292 N33292 0 diode
R33293 N33292 N33293 10
D33293 N33293 0 diode
R33294 N33293 N33294 10
D33294 N33294 0 diode
R33295 N33294 N33295 10
D33295 N33295 0 diode
R33296 N33295 N33296 10
D33296 N33296 0 diode
R33297 N33296 N33297 10
D33297 N33297 0 diode
R33298 N33297 N33298 10
D33298 N33298 0 diode
R33299 N33298 N33299 10
D33299 N33299 0 diode
R33300 N33299 N33300 10
D33300 N33300 0 diode
R33301 N33300 N33301 10
D33301 N33301 0 diode
R33302 N33301 N33302 10
D33302 N33302 0 diode
R33303 N33302 N33303 10
D33303 N33303 0 diode
R33304 N33303 N33304 10
D33304 N33304 0 diode
R33305 N33304 N33305 10
D33305 N33305 0 diode
R33306 N33305 N33306 10
D33306 N33306 0 diode
R33307 N33306 N33307 10
D33307 N33307 0 diode
R33308 N33307 N33308 10
D33308 N33308 0 diode
R33309 N33308 N33309 10
D33309 N33309 0 diode
R33310 N33309 N33310 10
D33310 N33310 0 diode
R33311 N33310 N33311 10
D33311 N33311 0 diode
R33312 N33311 N33312 10
D33312 N33312 0 diode
R33313 N33312 N33313 10
D33313 N33313 0 diode
R33314 N33313 N33314 10
D33314 N33314 0 diode
R33315 N33314 N33315 10
D33315 N33315 0 diode
R33316 N33315 N33316 10
D33316 N33316 0 diode
R33317 N33316 N33317 10
D33317 N33317 0 diode
R33318 N33317 N33318 10
D33318 N33318 0 diode
R33319 N33318 N33319 10
D33319 N33319 0 diode
R33320 N33319 N33320 10
D33320 N33320 0 diode
R33321 N33320 N33321 10
D33321 N33321 0 diode
R33322 N33321 N33322 10
D33322 N33322 0 diode
R33323 N33322 N33323 10
D33323 N33323 0 diode
R33324 N33323 N33324 10
D33324 N33324 0 diode
R33325 N33324 N33325 10
D33325 N33325 0 diode
R33326 N33325 N33326 10
D33326 N33326 0 diode
R33327 N33326 N33327 10
D33327 N33327 0 diode
R33328 N33327 N33328 10
D33328 N33328 0 diode
R33329 N33328 N33329 10
D33329 N33329 0 diode
R33330 N33329 N33330 10
D33330 N33330 0 diode
R33331 N33330 N33331 10
D33331 N33331 0 diode
R33332 N33331 N33332 10
D33332 N33332 0 diode
R33333 N33332 N33333 10
D33333 N33333 0 diode
R33334 N33333 N33334 10
D33334 N33334 0 diode
R33335 N33334 N33335 10
D33335 N33335 0 diode
R33336 N33335 N33336 10
D33336 N33336 0 diode
R33337 N33336 N33337 10
D33337 N33337 0 diode
R33338 N33337 N33338 10
D33338 N33338 0 diode
R33339 N33338 N33339 10
D33339 N33339 0 diode
R33340 N33339 N33340 10
D33340 N33340 0 diode
R33341 N33340 N33341 10
D33341 N33341 0 diode
R33342 N33341 N33342 10
D33342 N33342 0 diode
R33343 N33342 N33343 10
D33343 N33343 0 diode
R33344 N33343 N33344 10
D33344 N33344 0 diode
R33345 N33344 N33345 10
D33345 N33345 0 diode
R33346 N33345 N33346 10
D33346 N33346 0 diode
R33347 N33346 N33347 10
D33347 N33347 0 diode
R33348 N33347 N33348 10
D33348 N33348 0 diode
R33349 N33348 N33349 10
D33349 N33349 0 diode
R33350 N33349 N33350 10
D33350 N33350 0 diode
R33351 N33350 N33351 10
D33351 N33351 0 diode
R33352 N33351 N33352 10
D33352 N33352 0 diode
R33353 N33352 N33353 10
D33353 N33353 0 diode
R33354 N33353 N33354 10
D33354 N33354 0 diode
R33355 N33354 N33355 10
D33355 N33355 0 diode
R33356 N33355 N33356 10
D33356 N33356 0 diode
R33357 N33356 N33357 10
D33357 N33357 0 diode
R33358 N33357 N33358 10
D33358 N33358 0 diode
R33359 N33358 N33359 10
D33359 N33359 0 diode
R33360 N33359 N33360 10
D33360 N33360 0 diode
R33361 N33360 N33361 10
D33361 N33361 0 diode
R33362 N33361 N33362 10
D33362 N33362 0 diode
R33363 N33362 N33363 10
D33363 N33363 0 diode
R33364 N33363 N33364 10
D33364 N33364 0 diode
R33365 N33364 N33365 10
D33365 N33365 0 diode
R33366 N33365 N33366 10
D33366 N33366 0 diode
R33367 N33366 N33367 10
D33367 N33367 0 diode
R33368 N33367 N33368 10
D33368 N33368 0 diode
R33369 N33368 N33369 10
D33369 N33369 0 diode
R33370 N33369 N33370 10
D33370 N33370 0 diode
R33371 N33370 N33371 10
D33371 N33371 0 diode
R33372 N33371 N33372 10
D33372 N33372 0 diode
R33373 N33372 N33373 10
D33373 N33373 0 diode
R33374 N33373 N33374 10
D33374 N33374 0 diode
R33375 N33374 N33375 10
D33375 N33375 0 diode
R33376 N33375 N33376 10
D33376 N33376 0 diode
R33377 N33376 N33377 10
D33377 N33377 0 diode
R33378 N33377 N33378 10
D33378 N33378 0 diode
R33379 N33378 N33379 10
D33379 N33379 0 diode
R33380 N33379 N33380 10
D33380 N33380 0 diode
R33381 N33380 N33381 10
D33381 N33381 0 diode
R33382 N33381 N33382 10
D33382 N33382 0 diode
R33383 N33382 N33383 10
D33383 N33383 0 diode
R33384 N33383 N33384 10
D33384 N33384 0 diode
R33385 N33384 N33385 10
D33385 N33385 0 diode
R33386 N33385 N33386 10
D33386 N33386 0 diode
R33387 N33386 N33387 10
D33387 N33387 0 diode
R33388 N33387 N33388 10
D33388 N33388 0 diode
R33389 N33388 N33389 10
D33389 N33389 0 diode
R33390 N33389 N33390 10
D33390 N33390 0 diode
R33391 N33390 N33391 10
D33391 N33391 0 diode
R33392 N33391 N33392 10
D33392 N33392 0 diode
R33393 N33392 N33393 10
D33393 N33393 0 diode
R33394 N33393 N33394 10
D33394 N33394 0 diode
R33395 N33394 N33395 10
D33395 N33395 0 diode
R33396 N33395 N33396 10
D33396 N33396 0 diode
R33397 N33396 N33397 10
D33397 N33397 0 diode
R33398 N33397 N33398 10
D33398 N33398 0 diode
R33399 N33398 N33399 10
D33399 N33399 0 diode
R33400 N33399 N33400 10
D33400 N33400 0 diode
R33401 N33400 N33401 10
D33401 N33401 0 diode
R33402 N33401 N33402 10
D33402 N33402 0 diode
R33403 N33402 N33403 10
D33403 N33403 0 diode
R33404 N33403 N33404 10
D33404 N33404 0 diode
R33405 N33404 N33405 10
D33405 N33405 0 diode
R33406 N33405 N33406 10
D33406 N33406 0 diode
R33407 N33406 N33407 10
D33407 N33407 0 diode
R33408 N33407 N33408 10
D33408 N33408 0 diode
R33409 N33408 N33409 10
D33409 N33409 0 diode
R33410 N33409 N33410 10
D33410 N33410 0 diode
R33411 N33410 N33411 10
D33411 N33411 0 diode
R33412 N33411 N33412 10
D33412 N33412 0 diode
R33413 N33412 N33413 10
D33413 N33413 0 diode
R33414 N33413 N33414 10
D33414 N33414 0 diode
R33415 N33414 N33415 10
D33415 N33415 0 diode
R33416 N33415 N33416 10
D33416 N33416 0 diode
R33417 N33416 N33417 10
D33417 N33417 0 diode
R33418 N33417 N33418 10
D33418 N33418 0 diode
R33419 N33418 N33419 10
D33419 N33419 0 diode
R33420 N33419 N33420 10
D33420 N33420 0 diode
R33421 N33420 N33421 10
D33421 N33421 0 diode
R33422 N33421 N33422 10
D33422 N33422 0 diode
R33423 N33422 N33423 10
D33423 N33423 0 diode
R33424 N33423 N33424 10
D33424 N33424 0 diode
R33425 N33424 N33425 10
D33425 N33425 0 diode
R33426 N33425 N33426 10
D33426 N33426 0 diode
R33427 N33426 N33427 10
D33427 N33427 0 diode
R33428 N33427 N33428 10
D33428 N33428 0 diode
R33429 N33428 N33429 10
D33429 N33429 0 diode
R33430 N33429 N33430 10
D33430 N33430 0 diode
R33431 N33430 N33431 10
D33431 N33431 0 diode
R33432 N33431 N33432 10
D33432 N33432 0 diode
R33433 N33432 N33433 10
D33433 N33433 0 diode
R33434 N33433 N33434 10
D33434 N33434 0 diode
R33435 N33434 N33435 10
D33435 N33435 0 diode
R33436 N33435 N33436 10
D33436 N33436 0 diode
R33437 N33436 N33437 10
D33437 N33437 0 diode
R33438 N33437 N33438 10
D33438 N33438 0 diode
R33439 N33438 N33439 10
D33439 N33439 0 diode
R33440 N33439 N33440 10
D33440 N33440 0 diode
R33441 N33440 N33441 10
D33441 N33441 0 diode
R33442 N33441 N33442 10
D33442 N33442 0 diode
R33443 N33442 N33443 10
D33443 N33443 0 diode
R33444 N33443 N33444 10
D33444 N33444 0 diode
R33445 N33444 N33445 10
D33445 N33445 0 diode
R33446 N33445 N33446 10
D33446 N33446 0 diode
R33447 N33446 N33447 10
D33447 N33447 0 diode
R33448 N33447 N33448 10
D33448 N33448 0 diode
R33449 N33448 N33449 10
D33449 N33449 0 diode
R33450 N33449 N33450 10
D33450 N33450 0 diode
R33451 N33450 N33451 10
D33451 N33451 0 diode
R33452 N33451 N33452 10
D33452 N33452 0 diode
R33453 N33452 N33453 10
D33453 N33453 0 diode
R33454 N33453 N33454 10
D33454 N33454 0 diode
R33455 N33454 N33455 10
D33455 N33455 0 diode
R33456 N33455 N33456 10
D33456 N33456 0 diode
R33457 N33456 N33457 10
D33457 N33457 0 diode
R33458 N33457 N33458 10
D33458 N33458 0 diode
R33459 N33458 N33459 10
D33459 N33459 0 diode
R33460 N33459 N33460 10
D33460 N33460 0 diode
R33461 N33460 N33461 10
D33461 N33461 0 diode
R33462 N33461 N33462 10
D33462 N33462 0 diode
R33463 N33462 N33463 10
D33463 N33463 0 diode
R33464 N33463 N33464 10
D33464 N33464 0 diode
R33465 N33464 N33465 10
D33465 N33465 0 diode
R33466 N33465 N33466 10
D33466 N33466 0 diode
R33467 N33466 N33467 10
D33467 N33467 0 diode
R33468 N33467 N33468 10
D33468 N33468 0 diode
R33469 N33468 N33469 10
D33469 N33469 0 diode
R33470 N33469 N33470 10
D33470 N33470 0 diode
R33471 N33470 N33471 10
D33471 N33471 0 diode
R33472 N33471 N33472 10
D33472 N33472 0 diode
R33473 N33472 N33473 10
D33473 N33473 0 diode
R33474 N33473 N33474 10
D33474 N33474 0 diode
R33475 N33474 N33475 10
D33475 N33475 0 diode
R33476 N33475 N33476 10
D33476 N33476 0 diode
R33477 N33476 N33477 10
D33477 N33477 0 diode
R33478 N33477 N33478 10
D33478 N33478 0 diode
R33479 N33478 N33479 10
D33479 N33479 0 diode
R33480 N33479 N33480 10
D33480 N33480 0 diode
R33481 N33480 N33481 10
D33481 N33481 0 diode
R33482 N33481 N33482 10
D33482 N33482 0 diode
R33483 N33482 N33483 10
D33483 N33483 0 diode
R33484 N33483 N33484 10
D33484 N33484 0 diode
R33485 N33484 N33485 10
D33485 N33485 0 diode
R33486 N33485 N33486 10
D33486 N33486 0 diode
R33487 N33486 N33487 10
D33487 N33487 0 diode
R33488 N33487 N33488 10
D33488 N33488 0 diode
R33489 N33488 N33489 10
D33489 N33489 0 diode
R33490 N33489 N33490 10
D33490 N33490 0 diode
R33491 N33490 N33491 10
D33491 N33491 0 diode
R33492 N33491 N33492 10
D33492 N33492 0 diode
R33493 N33492 N33493 10
D33493 N33493 0 diode
R33494 N33493 N33494 10
D33494 N33494 0 diode
R33495 N33494 N33495 10
D33495 N33495 0 diode
R33496 N33495 N33496 10
D33496 N33496 0 diode
R33497 N33496 N33497 10
D33497 N33497 0 diode
R33498 N33497 N33498 10
D33498 N33498 0 diode
R33499 N33498 N33499 10
D33499 N33499 0 diode
R33500 N33499 N33500 10
D33500 N33500 0 diode
R33501 N33500 N33501 10
D33501 N33501 0 diode
R33502 N33501 N33502 10
D33502 N33502 0 diode
R33503 N33502 N33503 10
D33503 N33503 0 diode
R33504 N33503 N33504 10
D33504 N33504 0 diode
R33505 N33504 N33505 10
D33505 N33505 0 diode
R33506 N33505 N33506 10
D33506 N33506 0 diode
R33507 N33506 N33507 10
D33507 N33507 0 diode
R33508 N33507 N33508 10
D33508 N33508 0 diode
R33509 N33508 N33509 10
D33509 N33509 0 diode
R33510 N33509 N33510 10
D33510 N33510 0 diode
R33511 N33510 N33511 10
D33511 N33511 0 diode
R33512 N33511 N33512 10
D33512 N33512 0 diode
R33513 N33512 N33513 10
D33513 N33513 0 diode
R33514 N33513 N33514 10
D33514 N33514 0 diode
R33515 N33514 N33515 10
D33515 N33515 0 diode
R33516 N33515 N33516 10
D33516 N33516 0 diode
R33517 N33516 N33517 10
D33517 N33517 0 diode
R33518 N33517 N33518 10
D33518 N33518 0 diode
R33519 N33518 N33519 10
D33519 N33519 0 diode
R33520 N33519 N33520 10
D33520 N33520 0 diode
R33521 N33520 N33521 10
D33521 N33521 0 diode
R33522 N33521 N33522 10
D33522 N33522 0 diode
R33523 N33522 N33523 10
D33523 N33523 0 diode
R33524 N33523 N33524 10
D33524 N33524 0 diode
R33525 N33524 N33525 10
D33525 N33525 0 diode
R33526 N33525 N33526 10
D33526 N33526 0 diode
R33527 N33526 N33527 10
D33527 N33527 0 diode
R33528 N33527 N33528 10
D33528 N33528 0 diode
R33529 N33528 N33529 10
D33529 N33529 0 diode
R33530 N33529 N33530 10
D33530 N33530 0 diode
R33531 N33530 N33531 10
D33531 N33531 0 diode
R33532 N33531 N33532 10
D33532 N33532 0 diode
R33533 N33532 N33533 10
D33533 N33533 0 diode
R33534 N33533 N33534 10
D33534 N33534 0 diode
R33535 N33534 N33535 10
D33535 N33535 0 diode
R33536 N33535 N33536 10
D33536 N33536 0 diode
R33537 N33536 N33537 10
D33537 N33537 0 diode
R33538 N33537 N33538 10
D33538 N33538 0 diode
R33539 N33538 N33539 10
D33539 N33539 0 diode
R33540 N33539 N33540 10
D33540 N33540 0 diode
R33541 N33540 N33541 10
D33541 N33541 0 diode
R33542 N33541 N33542 10
D33542 N33542 0 diode
R33543 N33542 N33543 10
D33543 N33543 0 diode
R33544 N33543 N33544 10
D33544 N33544 0 diode
R33545 N33544 N33545 10
D33545 N33545 0 diode
R33546 N33545 N33546 10
D33546 N33546 0 diode
R33547 N33546 N33547 10
D33547 N33547 0 diode
R33548 N33547 N33548 10
D33548 N33548 0 diode
R33549 N33548 N33549 10
D33549 N33549 0 diode
R33550 N33549 N33550 10
D33550 N33550 0 diode
R33551 N33550 N33551 10
D33551 N33551 0 diode
R33552 N33551 N33552 10
D33552 N33552 0 diode
R33553 N33552 N33553 10
D33553 N33553 0 diode
R33554 N33553 N33554 10
D33554 N33554 0 diode
R33555 N33554 N33555 10
D33555 N33555 0 diode
R33556 N33555 N33556 10
D33556 N33556 0 diode
R33557 N33556 N33557 10
D33557 N33557 0 diode
R33558 N33557 N33558 10
D33558 N33558 0 diode
R33559 N33558 N33559 10
D33559 N33559 0 diode
R33560 N33559 N33560 10
D33560 N33560 0 diode
R33561 N33560 N33561 10
D33561 N33561 0 diode
R33562 N33561 N33562 10
D33562 N33562 0 diode
R33563 N33562 N33563 10
D33563 N33563 0 diode
R33564 N33563 N33564 10
D33564 N33564 0 diode
R33565 N33564 N33565 10
D33565 N33565 0 diode
R33566 N33565 N33566 10
D33566 N33566 0 diode
R33567 N33566 N33567 10
D33567 N33567 0 diode
R33568 N33567 N33568 10
D33568 N33568 0 diode
R33569 N33568 N33569 10
D33569 N33569 0 diode
R33570 N33569 N33570 10
D33570 N33570 0 diode
R33571 N33570 N33571 10
D33571 N33571 0 diode
R33572 N33571 N33572 10
D33572 N33572 0 diode
R33573 N33572 N33573 10
D33573 N33573 0 diode
R33574 N33573 N33574 10
D33574 N33574 0 diode
R33575 N33574 N33575 10
D33575 N33575 0 diode
R33576 N33575 N33576 10
D33576 N33576 0 diode
R33577 N33576 N33577 10
D33577 N33577 0 diode
R33578 N33577 N33578 10
D33578 N33578 0 diode
R33579 N33578 N33579 10
D33579 N33579 0 diode
R33580 N33579 N33580 10
D33580 N33580 0 diode
R33581 N33580 N33581 10
D33581 N33581 0 diode
R33582 N33581 N33582 10
D33582 N33582 0 diode
R33583 N33582 N33583 10
D33583 N33583 0 diode
R33584 N33583 N33584 10
D33584 N33584 0 diode
R33585 N33584 N33585 10
D33585 N33585 0 diode
R33586 N33585 N33586 10
D33586 N33586 0 diode
R33587 N33586 N33587 10
D33587 N33587 0 diode
R33588 N33587 N33588 10
D33588 N33588 0 diode
R33589 N33588 N33589 10
D33589 N33589 0 diode
R33590 N33589 N33590 10
D33590 N33590 0 diode
R33591 N33590 N33591 10
D33591 N33591 0 diode
R33592 N33591 N33592 10
D33592 N33592 0 diode
R33593 N33592 N33593 10
D33593 N33593 0 diode
R33594 N33593 N33594 10
D33594 N33594 0 diode
R33595 N33594 N33595 10
D33595 N33595 0 diode
R33596 N33595 N33596 10
D33596 N33596 0 diode
R33597 N33596 N33597 10
D33597 N33597 0 diode
R33598 N33597 N33598 10
D33598 N33598 0 diode
R33599 N33598 N33599 10
D33599 N33599 0 diode
R33600 N33599 N33600 10
D33600 N33600 0 diode
R33601 N33600 N33601 10
D33601 N33601 0 diode
R33602 N33601 N33602 10
D33602 N33602 0 diode
R33603 N33602 N33603 10
D33603 N33603 0 diode
R33604 N33603 N33604 10
D33604 N33604 0 diode
R33605 N33604 N33605 10
D33605 N33605 0 diode
R33606 N33605 N33606 10
D33606 N33606 0 diode
R33607 N33606 N33607 10
D33607 N33607 0 diode
R33608 N33607 N33608 10
D33608 N33608 0 diode
R33609 N33608 N33609 10
D33609 N33609 0 diode
R33610 N33609 N33610 10
D33610 N33610 0 diode
R33611 N33610 N33611 10
D33611 N33611 0 diode
R33612 N33611 N33612 10
D33612 N33612 0 diode
R33613 N33612 N33613 10
D33613 N33613 0 diode
R33614 N33613 N33614 10
D33614 N33614 0 diode
R33615 N33614 N33615 10
D33615 N33615 0 diode
R33616 N33615 N33616 10
D33616 N33616 0 diode
R33617 N33616 N33617 10
D33617 N33617 0 diode
R33618 N33617 N33618 10
D33618 N33618 0 diode
R33619 N33618 N33619 10
D33619 N33619 0 diode
R33620 N33619 N33620 10
D33620 N33620 0 diode
R33621 N33620 N33621 10
D33621 N33621 0 diode
R33622 N33621 N33622 10
D33622 N33622 0 diode
R33623 N33622 N33623 10
D33623 N33623 0 diode
R33624 N33623 N33624 10
D33624 N33624 0 diode
R33625 N33624 N33625 10
D33625 N33625 0 diode
R33626 N33625 N33626 10
D33626 N33626 0 diode
R33627 N33626 N33627 10
D33627 N33627 0 diode
R33628 N33627 N33628 10
D33628 N33628 0 diode
R33629 N33628 N33629 10
D33629 N33629 0 diode
R33630 N33629 N33630 10
D33630 N33630 0 diode
R33631 N33630 N33631 10
D33631 N33631 0 diode
R33632 N33631 N33632 10
D33632 N33632 0 diode
R33633 N33632 N33633 10
D33633 N33633 0 diode
R33634 N33633 N33634 10
D33634 N33634 0 diode
R33635 N33634 N33635 10
D33635 N33635 0 diode
R33636 N33635 N33636 10
D33636 N33636 0 diode
R33637 N33636 N33637 10
D33637 N33637 0 diode
R33638 N33637 N33638 10
D33638 N33638 0 diode
R33639 N33638 N33639 10
D33639 N33639 0 diode
R33640 N33639 N33640 10
D33640 N33640 0 diode
R33641 N33640 N33641 10
D33641 N33641 0 diode
R33642 N33641 N33642 10
D33642 N33642 0 diode
R33643 N33642 N33643 10
D33643 N33643 0 diode
R33644 N33643 N33644 10
D33644 N33644 0 diode
R33645 N33644 N33645 10
D33645 N33645 0 diode
R33646 N33645 N33646 10
D33646 N33646 0 diode
R33647 N33646 N33647 10
D33647 N33647 0 diode
R33648 N33647 N33648 10
D33648 N33648 0 diode
R33649 N33648 N33649 10
D33649 N33649 0 diode
R33650 N33649 N33650 10
D33650 N33650 0 diode
R33651 N33650 N33651 10
D33651 N33651 0 diode
R33652 N33651 N33652 10
D33652 N33652 0 diode
R33653 N33652 N33653 10
D33653 N33653 0 diode
R33654 N33653 N33654 10
D33654 N33654 0 diode
R33655 N33654 N33655 10
D33655 N33655 0 diode
R33656 N33655 N33656 10
D33656 N33656 0 diode
R33657 N33656 N33657 10
D33657 N33657 0 diode
R33658 N33657 N33658 10
D33658 N33658 0 diode
R33659 N33658 N33659 10
D33659 N33659 0 diode
R33660 N33659 N33660 10
D33660 N33660 0 diode
R33661 N33660 N33661 10
D33661 N33661 0 diode
R33662 N33661 N33662 10
D33662 N33662 0 diode
R33663 N33662 N33663 10
D33663 N33663 0 diode
R33664 N33663 N33664 10
D33664 N33664 0 diode
R33665 N33664 N33665 10
D33665 N33665 0 diode
R33666 N33665 N33666 10
D33666 N33666 0 diode
R33667 N33666 N33667 10
D33667 N33667 0 diode
R33668 N33667 N33668 10
D33668 N33668 0 diode
R33669 N33668 N33669 10
D33669 N33669 0 diode
R33670 N33669 N33670 10
D33670 N33670 0 diode
R33671 N33670 N33671 10
D33671 N33671 0 diode
R33672 N33671 N33672 10
D33672 N33672 0 diode
R33673 N33672 N33673 10
D33673 N33673 0 diode
R33674 N33673 N33674 10
D33674 N33674 0 diode
R33675 N33674 N33675 10
D33675 N33675 0 diode
R33676 N33675 N33676 10
D33676 N33676 0 diode
R33677 N33676 N33677 10
D33677 N33677 0 diode
R33678 N33677 N33678 10
D33678 N33678 0 diode
R33679 N33678 N33679 10
D33679 N33679 0 diode
R33680 N33679 N33680 10
D33680 N33680 0 diode
R33681 N33680 N33681 10
D33681 N33681 0 diode
R33682 N33681 N33682 10
D33682 N33682 0 diode
R33683 N33682 N33683 10
D33683 N33683 0 diode
R33684 N33683 N33684 10
D33684 N33684 0 diode
R33685 N33684 N33685 10
D33685 N33685 0 diode
R33686 N33685 N33686 10
D33686 N33686 0 diode
R33687 N33686 N33687 10
D33687 N33687 0 diode
R33688 N33687 N33688 10
D33688 N33688 0 diode
R33689 N33688 N33689 10
D33689 N33689 0 diode
R33690 N33689 N33690 10
D33690 N33690 0 diode
R33691 N33690 N33691 10
D33691 N33691 0 diode
R33692 N33691 N33692 10
D33692 N33692 0 diode
R33693 N33692 N33693 10
D33693 N33693 0 diode
R33694 N33693 N33694 10
D33694 N33694 0 diode
R33695 N33694 N33695 10
D33695 N33695 0 diode
R33696 N33695 N33696 10
D33696 N33696 0 diode
R33697 N33696 N33697 10
D33697 N33697 0 diode
R33698 N33697 N33698 10
D33698 N33698 0 diode
R33699 N33698 N33699 10
D33699 N33699 0 diode
R33700 N33699 N33700 10
D33700 N33700 0 diode
R33701 N33700 N33701 10
D33701 N33701 0 diode
R33702 N33701 N33702 10
D33702 N33702 0 diode
R33703 N33702 N33703 10
D33703 N33703 0 diode
R33704 N33703 N33704 10
D33704 N33704 0 diode
R33705 N33704 N33705 10
D33705 N33705 0 diode
R33706 N33705 N33706 10
D33706 N33706 0 diode
R33707 N33706 N33707 10
D33707 N33707 0 diode
R33708 N33707 N33708 10
D33708 N33708 0 diode
R33709 N33708 N33709 10
D33709 N33709 0 diode
R33710 N33709 N33710 10
D33710 N33710 0 diode
R33711 N33710 N33711 10
D33711 N33711 0 diode
R33712 N33711 N33712 10
D33712 N33712 0 diode
R33713 N33712 N33713 10
D33713 N33713 0 diode
R33714 N33713 N33714 10
D33714 N33714 0 diode
R33715 N33714 N33715 10
D33715 N33715 0 diode
R33716 N33715 N33716 10
D33716 N33716 0 diode
R33717 N33716 N33717 10
D33717 N33717 0 diode
R33718 N33717 N33718 10
D33718 N33718 0 diode
R33719 N33718 N33719 10
D33719 N33719 0 diode
R33720 N33719 N33720 10
D33720 N33720 0 diode
R33721 N33720 N33721 10
D33721 N33721 0 diode
R33722 N33721 N33722 10
D33722 N33722 0 diode
R33723 N33722 N33723 10
D33723 N33723 0 diode
R33724 N33723 N33724 10
D33724 N33724 0 diode
R33725 N33724 N33725 10
D33725 N33725 0 diode
R33726 N33725 N33726 10
D33726 N33726 0 diode
R33727 N33726 N33727 10
D33727 N33727 0 diode
R33728 N33727 N33728 10
D33728 N33728 0 diode
R33729 N33728 N33729 10
D33729 N33729 0 diode
R33730 N33729 N33730 10
D33730 N33730 0 diode
R33731 N33730 N33731 10
D33731 N33731 0 diode
R33732 N33731 N33732 10
D33732 N33732 0 diode
R33733 N33732 N33733 10
D33733 N33733 0 diode
R33734 N33733 N33734 10
D33734 N33734 0 diode
R33735 N33734 N33735 10
D33735 N33735 0 diode
R33736 N33735 N33736 10
D33736 N33736 0 diode
R33737 N33736 N33737 10
D33737 N33737 0 diode
R33738 N33737 N33738 10
D33738 N33738 0 diode
R33739 N33738 N33739 10
D33739 N33739 0 diode
R33740 N33739 N33740 10
D33740 N33740 0 diode
R33741 N33740 N33741 10
D33741 N33741 0 diode
R33742 N33741 N33742 10
D33742 N33742 0 diode
R33743 N33742 N33743 10
D33743 N33743 0 diode
R33744 N33743 N33744 10
D33744 N33744 0 diode
R33745 N33744 N33745 10
D33745 N33745 0 diode
R33746 N33745 N33746 10
D33746 N33746 0 diode
R33747 N33746 N33747 10
D33747 N33747 0 diode
R33748 N33747 N33748 10
D33748 N33748 0 diode
R33749 N33748 N33749 10
D33749 N33749 0 diode
R33750 N33749 N33750 10
D33750 N33750 0 diode
R33751 N33750 N33751 10
D33751 N33751 0 diode
R33752 N33751 N33752 10
D33752 N33752 0 diode
R33753 N33752 N33753 10
D33753 N33753 0 diode
R33754 N33753 N33754 10
D33754 N33754 0 diode
R33755 N33754 N33755 10
D33755 N33755 0 diode
R33756 N33755 N33756 10
D33756 N33756 0 diode
R33757 N33756 N33757 10
D33757 N33757 0 diode
R33758 N33757 N33758 10
D33758 N33758 0 diode
R33759 N33758 N33759 10
D33759 N33759 0 diode
R33760 N33759 N33760 10
D33760 N33760 0 diode
R33761 N33760 N33761 10
D33761 N33761 0 diode
R33762 N33761 N33762 10
D33762 N33762 0 diode
R33763 N33762 N33763 10
D33763 N33763 0 diode
R33764 N33763 N33764 10
D33764 N33764 0 diode
R33765 N33764 N33765 10
D33765 N33765 0 diode
R33766 N33765 N33766 10
D33766 N33766 0 diode
R33767 N33766 N33767 10
D33767 N33767 0 diode
R33768 N33767 N33768 10
D33768 N33768 0 diode
R33769 N33768 N33769 10
D33769 N33769 0 diode
R33770 N33769 N33770 10
D33770 N33770 0 diode
R33771 N33770 N33771 10
D33771 N33771 0 diode
R33772 N33771 N33772 10
D33772 N33772 0 diode
R33773 N33772 N33773 10
D33773 N33773 0 diode
R33774 N33773 N33774 10
D33774 N33774 0 diode
R33775 N33774 N33775 10
D33775 N33775 0 diode
R33776 N33775 N33776 10
D33776 N33776 0 diode
R33777 N33776 N33777 10
D33777 N33777 0 diode
R33778 N33777 N33778 10
D33778 N33778 0 diode
R33779 N33778 N33779 10
D33779 N33779 0 diode
R33780 N33779 N33780 10
D33780 N33780 0 diode
R33781 N33780 N33781 10
D33781 N33781 0 diode
R33782 N33781 N33782 10
D33782 N33782 0 diode
R33783 N33782 N33783 10
D33783 N33783 0 diode
R33784 N33783 N33784 10
D33784 N33784 0 diode
R33785 N33784 N33785 10
D33785 N33785 0 diode
R33786 N33785 N33786 10
D33786 N33786 0 diode
R33787 N33786 N33787 10
D33787 N33787 0 diode
R33788 N33787 N33788 10
D33788 N33788 0 diode
R33789 N33788 N33789 10
D33789 N33789 0 diode
R33790 N33789 N33790 10
D33790 N33790 0 diode
R33791 N33790 N33791 10
D33791 N33791 0 diode
R33792 N33791 N33792 10
D33792 N33792 0 diode
R33793 N33792 N33793 10
D33793 N33793 0 diode
R33794 N33793 N33794 10
D33794 N33794 0 diode
R33795 N33794 N33795 10
D33795 N33795 0 diode
R33796 N33795 N33796 10
D33796 N33796 0 diode
R33797 N33796 N33797 10
D33797 N33797 0 diode
R33798 N33797 N33798 10
D33798 N33798 0 diode
R33799 N33798 N33799 10
D33799 N33799 0 diode
R33800 N33799 N33800 10
D33800 N33800 0 diode
R33801 N33800 N33801 10
D33801 N33801 0 diode
R33802 N33801 N33802 10
D33802 N33802 0 diode
R33803 N33802 N33803 10
D33803 N33803 0 diode
R33804 N33803 N33804 10
D33804 N33804 0 diode
R33805 N33804 N33805 10
D33805 N33805 0 diode
R33806 N33805 N33806 10
D33806 N33806 0 diode
R33807 N33806 N33807 10
D33807 N33807 0 diode
R33808 N33807 N33808 10
D33808 N33808 0 diode
R33809 N33808 N33809 10
D33809 N33809 0 diode
R33810 N33809 N33810 10
D33810 N33810 0 diode
R33811 N33810 N33811 10
D33811 N33811 0 diode
R33812 N33811 N33812 10
D33812 N33812 0 diode
R33813 N33812 N33813 10
D33813 N33813 0 diode
R33814 N33813 N33814 10
D33814 N33814 0 diode
R33815 N33814 N33815 10
D33815 N33815 0 diode
R33816 N33815 N33816 10
D33816 N33816 0 diode
R33817 N33816 N33817 10
D33817 N33817 0 diode
R33818 N33817 N33818 10
D33818 N33818 0 diode
R33819 N33818 N33819 10
D33819 N33819 0 diode
R33820 N33819 N33820 10
D33820 N33820 0 diode
R33821 N33820 N33821 10
D33821 N33821 0 diode
R33822 N33821 N33822 10
D33822 N33822 0 diode
R33823 N33822 N33823 10
D33823 N33823 0 diode
R33824 N33823 N33824 10
D33824 N33824 0 diode
R33825 N33824 N33825 10
D33825 N33825 0 diode
R33826 N33825 N33826 10
D33826 N33826 0 diode
R33827 N33826 N33827 10
D33827 N33827 0 diode
R33828 N33827 N33828 10
D33828 N33828 0 diode
R33829 N33828 N33829 10
D33829 N33829 0 diode
R33830 N33829 N33830 10
D33830 N33830 0 diode
R33831 N33830 N33831 10
D33831 N33831 0 diode
R33832 N33831 N33832 10
D33832 N33832 0 diode
R33833 N33832 N33833 10
D33833 N33833 0 diode
R33834 N33833 N33834 10
D33834 N33834 0 diode
R33835 N33834 N33835 10
D33835 N33835 0 diode
R33836 N33835 N33836 10
D33836 N33836 0 diode
R33837 N33836 N33837 10
D33837 N33837 0 diode
R33838 N33837 N33838 10
D33838 N33838 0 diode
R33839 N33838 N33839 10
D33839 N33839 0 diode
R33840 N33839 N33840 10
D33840 N33840 0 diode
R33841 N33840 N33841 10
D33841 N33841 0 diode
R33842 N33841 N33842 10
D33842 N33842 0 diode
R33843 N33842 N33843 10
D33843 N33843 0 diode
R33844 N33843 N33844 10
D33844 N33844 0 diode
R33845 N33844 N33845 10
D33845 N33845 0 diode
R33846 N33845 N33846 10
D33846 N33846 0 diode
R33847 N33846 N33847 10
D33847 N33847 0 diode
R33848 N33847 N33848 10
D33848 N33848 0 diode
R33849 N33848 N33849 10
D33849 N33849 0 diode
R33850 N33849 N33850 10
D33850 N33850 0 diode
R33851 N33850 N33851 10
D33851 N33851 0 diode
R33852 N33851 N33852 10
D33852 N33852 0 diode
R33853 N33852 N33853 10
D33853 N33853 0 diode
R33854 N33853 N33854 10
D33854 N33854 0 diode
R33855 N33854 N33855 10
D33855 N33855 0 diode
R33856 N33855 N33856 10
D33856 N33856 0 diode
R33857 N33856 N33857 10
D33857 N33857 0 diode
R33858 N33857 N33858 10
D33858 N33858 0 diode
R33859 N33858 N33859 10
D33859 N33859 0 diode
R33860 N33859 N33860 10
D33860 N33860 0 diode
R33861 N33860 N33861 10
D33861 N33861 0 diode
R33862 N33861 N33862 10
D33862 N33862 0 diode
R33863 N33862 N33863 10
D33863 N33863 0 diode
R33864 N33863 N33864 10
D33864 N33864 0 diode
R33865 N33864 N33865 10
D33865 N33865 0 diode
R33866 N33865 N33866 10
D33866 N33866 0 diode
R33867 N33866 N33867 10
D33867 N33867 0 diode
R33868 N33867 N33868 10
D33868 N33868 0 diode
R33869 N33868 N33869 10
D33869 N33869 0 diode
R33870 N33869 N33870 10
D33870 N33870 0 diode
R33871 N33870 N33871 10
D33871 N33871 0 diode
R33872 N33871 N33872 10
D33872 N33872 0 diode
R33873 N33872 N33873 10
D33873 N33873 0 diode
R33874 N33873 N33874 10
D33874 N33874 0 diode
R33875 N33874 N33875 10
D33875 N33875 0 diode
R33876 N33875 N33876 10
D33876 N33876 0 diode
R33877 N33876 N33877 10
D33877 N33877 0 diode
R33878 N33877 N33878 10
D33878 N33878 0 diode
R33879 N33878 N33879 10
D33879 N33879 0 diode
R33880 N33879 N33880 10
D33880 N33880 0 diode
R33881 N33880 N33881 10
D33881 N33881 0 diode
R33882 N33881 N33882 10
D33882 N33882 0 diode
R33883 N33882 N33883 10
D33883 N33883 0 diode
R33884 N33883 N33884 10
D33884 N33884 0 diode
R33885 N33884 N33885 10
D33885 N33885 0 diode
R33886 N33885 N33886 10
D33886 N33886 0 diode
R33887 N33886 N33887 10
D33887 N33887 0 diode
R33888 N33887 N33888 10
D33888 N33888 0 diode
R33889 N33888 N33889 10
D33889 N33889 0 diode
R33890 N33889 N33890 10
D33890 N33890 0 diode
R33891 N33890 N33891 10
D33891 N33891 0 diode
R33892 N33891 N33892 10
D33892 N33892 0 diode
R33893 N33892 N33893 10
D33893 N33893 0 diode
R33894 N33893 N33894 10
D33894 N33894 0 diode
R33895 N33894 N33895 10
D33895 N33895 0 diode
R33896 N33895 N33896 10
D33896 N33896 0 diode
R33897 N33896 N33897 10
D33897 N33897 0 diode
R33898 N33897 N33898 10
D33898 N33898 0 diode
R33899 N33898 N33899 10
D33899 N33899 0 diode
R33900 N33899 N33900 10
D33900 N33900 0 diode
R33901 N33900 N33901 10
D33901 N33901 0 diode
R33902 N33901 N33902 10
D33902 N33902 0 diode
R33903 N33902 N33903 10
D33903 N33903 0 diode
R33904 N33903 N33904 10
D33904 N33904 0 diode
R33905 N33904 N33905 10
D33905 N33905 0 diode
R33906 N33905 N33906 10
D33906 N33906 0 diode
R33907 N33906 N33907 10
D33907 N33907 0 diode
R33908 N33907 N33908 10
D33908 N33908 0 diode
R33909 N33908 N33909 10
D33909 N33909 0 diode
R33910 N33909 N33910 10
D33910 N33910 0 diode
R33911 N33910 N33911 10
D33911 N33911 0 diode
R33912 N33911 N33912 10
D33912 N33912 0 diode
R33913 N33912 N33913 10
D33913 N33913 0 diode
R33914 N33913 N33914 10
D33914 N33914 0 diode
R33915 N33914 N33915 10
D33915 N33915 0 diode
R33916 N33915 N33916 10
D33916 N33916 0 diode
R33917 N33916 N33917 10
D33917 N33917 0 diode
R33918 N33917 N33918 10
D33918 N33918 0 diode
R33919 N33918 N33919 10
D33919 N33919 0 diode
R33920 N33919 N33920 10
D33920 N33920 0 diode
R33921 N33920 N33921 10
D33921 N33921 0 diode
R33922 N33921 N33922 10
D33922 N33922 0 diode
R33923 N33922 N33923 10
D33923 N33923 0 diode
R33924 N33923 N33924 10
D33924 N33924 0 diode
R33925 N33924 N33925 10
D33925 N33925 0 diode
R33926 N33925 N33926 10
D33926 N33926 0 diode
R33927 N33926 N33927 10
D33927 N33927 0 diode
R33928 N33927 N33928 10
D33928 N33928 0 diode
R33929 N33928 N33929 10
D33929 N33929 0 diode
R33930 N33929 N33930 10
D33930 N33930 0 diode
R33931 N33930 N33931 10
D33931 N33931 0 diode
R33932 N33931 N33932 10
D33932 N33932 0 diode
R33933 N33932 N33933 10
D33933 N33933 0 diode
R33934 N33933 N33934 10
D33934 N33934 0 diode
R33935 N33934 N33935 10
D33935 N33935 0 diode
R33936 N33935 N33936 10
D33936 N33936 0 diode
R33937 N33936 N33937 10
D33937 N33937 0 diode
R33938 N33937 N33938 10
D33938 N33938 0 diode
R33939 N33938 N33939 10
D33939 N33939 0 diode
R33940 N33939 N33940 10
D33940 N33940 0 diode
R33941 N33940 N33941 10
D33941 N33941 0 diode
R33942 N33941 N33942 10
D33942 N33942 0 diode
R33943 N33942 N33943 10
D33943 N33943 0 diode
R33944 N33943 N33944 10
D33944 N33944 0 diode
R33945 N33944 N33945 10
D33945 N33945 0 diode
R33946 N33945 N33946 10
D33946 N33946 0 diode
R33947 N33946 N33947 10
D33947 N33947 0 diode
R33948 N33947 N33948 10
D33948 N33948 0 diode
R33949 N33948 N33949 10
D33949 N33949 0 diode
R33950 N33949 N33950 10
D33950 N33950 0 diode
R33951 N33950 N33951 10
D33951 N33951 0 diode
R33952 N33951 N33952 10
D33952 N33952 0 diode
R33953 N33952 N33953 10
D33953 N33953 0 diode
R33954 N33953 N33954 10
D33954 N33954 0 diode
R33955 N33954 N33955 10
D33955 N33955 0 diode
R33956 N33955 N33956 10
D33956 N33956 0 diode
R33957 N33956 N33957 10
D33957 N33957 0 diode
R33958 N33957 N33958 10
D33958 N33958 0 diode
R33959 N33958 N33959 10
D33959 N33959 0 diode
R33960 N33959 N33960 10
D33960 N33960 0 diode
R33961 N33960 N33961 10
D33961 N33961 0 diode
R33962 N33961 N33962 10
D33962 N33962 0 diode
R33963 N33962 N33963 10
D33963 N33963 0 diode
R33964 N33963 N33964 10
D33964 N33964 0 diode
R33965 N33964 N33965 10
D33965 N33965 0 diode
R33966 N33965 N33966 10
D33966 N33966 0 diode
R33967 N33966 N33967 10
D33967 N33967 0 diode
R33968 N33967 N33968 10
D33968 N33968 0 diode
R33969 N33968 N33969 10
D33969 N33969 0 diode
R33970 N33969 N33970 10
D33970 N33970 0 diode
R33971 N33970 N33971 10
D33971 N33971 0 diode
R33972 N33971 N33972 10
D33972 N33972 0 diode
R33973 N33972 N33973 10
D33973 N33973 0 diode
R33974 N33973 N33974 10
D33974 N33974 0 diode
R33975 N33974 N33975 10
D33975 N33975 0 diode
R33976 N33975 N33976 10
D33976 N33976 0 diode
R33977 N33976 N33977 10
D33977 N33977 0 diode
R33978 N33977 N33978 10
D33978 N33978 0 diode
R33979 N33978 N33979 10
D33979 N33979 0 diode
R33980 N33979 N33980 10
D33980 N33980 0 diode
R33981 N33980 N33981 10
D33981 N33981 0 diode
R33982 N33981 N33982 10
D33982 N33982 0 diode
R33983 N33982 N33983 10
D33983 N33983 0 diode
R33984 N33983 N33984 10
D33984 N33984 0 diode
R33985 N33984 N33985 10
D33985 N33985 0 diode
R33986 N33985 N33986 10
D33986 N33986 0 diode
R33987 N33986 N33987 10
D33987 N33987 0 diode
R33988 N33987 N33988 10
D33988 N33988 0 diode
R33989 N33988 N33989 10
D33989 N33989 0 diode
R33990 N33989 N33990 10
D33990 N33990 0 diode
R33991 N33990 N33991 10
D33991 N33991 0 diode
R33992 N33991 N33992 10
D33992 N33992 0 diode
R33993 N33992 N33993 10
D33993 N33993 0 diode
R33994 N33993 N33994 10
D33994 N33994 0 diode
R33995 N33994 N33995 10
D33995 N33995 0 diode
R33996 N33995 N33996 10
D33996 N33996 0 diode
R33997 N33996 N33997 10
D33997 N33997 0 diode
R33998 N33997 N33998 10
D33998 N33998 0 diode
R33999 N33998 N33999 10
D33999 N33999 0 diode
R34000 N33999 N34000 10
D34000 N34000 0 diode
R34001 N34000 N34001 10
D34001 N34001 0 diode
R34002 N34001 N34002 10
D34002 N34002 0 diode
R34003 N34002 N34003 10
D34003 N34003 0 diode
R34004 N34003 N34004 10
D34004 N34004 0 diode
R34005 N34004 N34005 10
D34005 N34005 0 diode
R34006 N34005 N34006 10
D34006 N34006 0 diode
R34007 N34006 N34007 10
D34007 N34007 0 diode
R34008 N34007 N34008 10
D34008 N34008 0 diode
R34009 N34008 N34009 10
D34009 N34009 0 diode
R34010 N34009 N34010 10
D34010 N34010 0 diode
R34011 N34010 N34011 10
D34011 N34011 0 diode
R34012 N34011 N34012 10
D34012 N34012 0 diode
R34013 N34012 N34013 10
D34013 N34013 0 diode
R34014 N34013 N34014 10
D34014 N34014 0 diode
R34015 N34014 N34015 10
D34015 N34015 0 diode
R34016 N34015 N34016 10
D34016 N34016 0 diode
R34017 N34016 N34017 10
D34017 N34017 0 diode
R34018 N34017 N34018 10
D34018 N34018 0 diode
R34019 N34018 N34019 10
D34019 N34019 0 diode
R34020 N34019 N34020 10
D34020 N34020 0 diode
R34021 N34020 N34021 10
D34021 N34021 0 diode
R34022 N34021 N34022 10
D34022 N34022 0 diode
R34023 N34022 N34023 10
D34023 N34023 0 diode
R34024 N34023 N34024 10
D34024 N34024 0 diode
R34025 N34024 N34025 10
D34025 N34025 0 diode
R34026 N34025 N34026 10
D34026 N34026 0 diode
R34027 N34026 N34027 10
D34027 N34027 0 diode
R34028 N34027 N34028 10
D34028 N34028 0 diode
R34029 N34028 N34029 10
D34029 N34029 0 diode
R34030 N34029 N34030 10
D34030 N34030 0 diode
R34031 N34030 N34031 10
D34031 N34031 0 diode
R34032 N34031 N34032 10
D34032 N34032 0 diode
R34033 N34032 N34033 10
D34033 N34033 0 diode
R34034 N34033 N34034 10
D34034 N34034 0 diode
R34035 N34034 N34035 10
D34035 N34035 0 diode
R34036 N34035 N34036 10
D34036 N34036 0 diode
R34037 N34036 N34037 10
D34037 N34037 0 diode
R34038 N34037 N34038 10
D34038 N34038 0 diode
R34039 N34038 N34039 10
D34039 N34039 0 diode
R34040 N34039 N34040 10
D34040 N34040 0 diode
R34041 N34040 N34041 10
D34041 N34041 0 diode
R34042 N34041 N34042 10
D34042 N34042 0 diode
R34043 N34042 N34043 10
D34043 N34043 0 diode
R34044 N34043 N34044 10
D34044 N34044 0 diode
R34045 N34044 N34045 10
D34045 N34045 0 diode
R34046 N34045 N34046 10
D34046 N34046 0 diode
R34047 N34046 N34047 10
D34047 N34047 0 diode
R34048 N34047 N34048 10
D34048 N34048 0 diode
R34049 N34048 N34049 10
D34049 N34049 0 diode
R34050 N34049 N34050 10
D34050 N34050 0 diode
R34051 N34050 N34051 10
D34051 N34051 0 diode
R34052 N34051 N34052 10
D34052 N34052 0 diode
R34053 N34052 N34053 10
D34053 N34053 0 diode
R34054 N34053 N34054 10
D34054 N34054 0 diode
R34055 N34054 N34055 10
D34055 N34055 0 diode
R34056 N34055 N34056 10
D34056 N34056 0 diode
R34057 N34056 N34057 10
D34057 N34057 0 diode
R34058 N34057 N34058 10
D34058 N34058 0 diode
R34059 N34058 N34059 10
D34059 N34059 0 diode
R34060 N34059 N34060 10
D34060 N34060 0 diode
R34061 N34060 N34061 10
D34061 N34061 0 diode
R34062 N34061 N34062 10
D34062 N34062 0 diode
R34063 N34062 N34063 10
D34063 N34063 0 diode
R34064 N34063 N34064 10
D34064 N34064 0 diode
R34065 N34064 N34065 10
D34065 N34065 0 diode
R34066 N34065 N34066 10
D34066 N34066 0 diode
R34067 N34066 N34067 10
D34067 N34067 0 diode
R34068 N34067 N34068 10
D34068 N34068 0 diode
R34069 N34068 N34069 10
D34069 N34069 0 diode
R34070 N34069 N34070 10
D34070 N34070 0 diode
R34071 N34070 N34071 10
D34071 N34071 0 diode
R34072 N34071 N34072 10
D34072 N34072 0 diode
R34073 N34072 N34073 10
D34073 N34073 0 diode
R34074 N34073 N34074 10
D34074 N34074 0 diode
R34075 N34074 N34075 10
D34075 N34075 0 diode
R34076 N34075 N34076 10
D34076 N34076 0 diode
R34077 N34076 N34077 10
D34077 N34077 0 diode
R34078 N34077 N34078 10
D34078 N34078 0 diode
R34079 N34078 N34079 10
D34079 N34079 0 diode
R34080 N34079 N34080 10
D34080 N34080 0 diode
R34081 N34080 N34081 10
D34081 N34081 0 diode
R34082 N34081 N34082 10
D34082 N34082 0 diode
R34083 N34082 N34083 10
D34083 N34083 0 diode
R34084 N34083 N34084 10
D34084 N34084 0 diode
R34085 N34084 N34085 10
D34085 N34085 0 diode
R34086 N34085 N34086 10
D34086 N34086 0 diode
R34087 N34086 N34087 10
D34087 N34087 0 diode
R34088 N34087 N34088 10
D34088 N34088 0 diode
R34089 N34088 N34089 10
D34089 N34089 0 diode
R34090 N34089 N34090 10
D34090 N34090 0 diode
R34091 N34090 N34091 10
D34091 N34091 0 diode
R34092 N34091 N34092 10
D34092 N34092 0 diode
R34093 N34092 N34093 10
D34093 N34093 0 diode
R34094 N34093 N34094 10
D34094 N34094 0 diode
R34095 N34094 N34095 10
D34095 N34095 0 diode
R34096 N34095 N34096 10
D34096 N34096 0 diode
R34097 N34096 N34097 10
D34097 N34097 0 diode
R34098 N34097 N34098 10
D34098 N34098 0 diode
R34099 N34098 N34099 10
D34099 N34099 0 diode
R34100 N34099 N34100 10
D34100 N34100 0 diode
R34101 N34100 N34101 10
D34101 N34101 0 diode
R34102 N34101 N34102 10
D34102 N34102 0 diode
R34103 N34102 N34103 10
D34103 N34103 0 diode
R34104 N34103 N34104 10
D34104 N34104 0 diode
R34105 N34104 N34105 10
D34105 N34105 0 diode
R34106 N34105 N34106 10
D34106 N34106 0 diode
R34107 N34106 N34107 10
D34107 N34107 0 diode
R34108 N34107 N34108 10
D34108 N34108 0 diode
R34109 N34108 N34109 10
D34109 N34109 0 diode
R34110 N34109 N34110 10
D34110 N34110 0 diode
R34111 N34110 N34111 10
D34111 N34111 0 diode
R34112 N34111 N34112 10
D34112 N34112 0 diode
R34113 N34112 N34113 10
D34113 N34113 0 diode
R34114 N34113 N34114 10
D34114 N34114 0 diode
R34115 N34114 N34115 10
D34115 N34115 0 diode
R34116 N34115 N34116 10
D34116 N34116 0 diode
R34117 N34116 N34117 10
D34117 N34117 0 diode
R34118 N34117 N34118 10
D34118 N34118 0 diode
R34119 N34118 N34119 10
D34119 N34119 0 diode
R34120 N34119 N34120 10
D34120 N34120 0 diode
R34121 N34120 N34121 10
D34121 N34121 0 diode
R34122 N34121 N34122 10
D34122 N34122 0 diode
R34123 N34122 N34123 10
D34123 N34123 0 diode
R34124 N34123 N34124 10
D34124 N34124 0 diode
R34125 N34124 N34125 10
D34125 N34125 0 diode
R34126 N34125 N34126 10
D34126 N34126 0 diode
R34127 N34126 N34127 10
D34127 N34127 0 diode
R34128 N34127 N34128 10
D34128 N34128 0 diode
R34129 N34128 N34129 10
D34129 N34129 0 diode
R34130 N34129 N34130 10
D34130 N34130 0 diode
R34131 N34130 N34131 10
D34131 N34131 0 diode
R34132 N34131 N34132 10
D34132 N34132 0 diode
R34133 N34132 N34133 10
D34133 N34133 0 diode
R34134 N34133 N34134 10
D34134 N34134 0 diode
R34135 N34134 N34135 10
D34135 N34135 0 diode
R34136 N34135 N34136 10
D34136 N34136 0 diode
R34137 N34136 N34137 10
D34137 N34137 0 diode
R34138 N34137 N34138 10
D34138 N34138 0 diode
R34139 N34138 N34139 10
D34139 N34139 0 diode
R34140 N34139 N34140 10
D34140 N34140 0 diode
R34141 N34140 N34141 10
D34141 N34141 0 diode
R34142 N34141 N34142 10
D34142 N34142 0 diode
R34143 N34142 N34143 10
D34143 N34143 0 diode
R34144 N34143 N34144 10
D34144 N34144 0 diode
R34145 N34144 N34145 10
D34145 N34145 0 diode
R34146 N34145 N34146 10
D34146 N34146 0 diode
R34147 N34146 N34147 10
D34147 N34147 0 diode
R34148 N34147 N34148 10
D34148 N34148 0 diode
R34149 N34148 N34149 10
D34149 N34149 0 diode
R34150 N34149 N34150 10
D34150 N34150 0 diode
R34151 N34150 N34151 10
D34151 N34151 0 diode
R34152 N34151 N34152 10
D34152 N34152 0 diode
R34153 N34152 N34153 10
D34153 N34153 0 diode
R34154 N34153 N34154 10
D34154 N34154 0 diode
R34155 N34154 N34155 10
D34155 N34155 0 diode
R34156 N34155 N34156 10
D34156 N34156 0 diode
R34157 N34156 N34157 10
D34157 N34157 0 diode
R34158 N34157 N34158 10
D34158 N34158 0 diode
R34159 N34158 N34159 10
D34159 N34159 0 diode
R34160 N34159 N34160 10
D34160 N34160 0 diode
R34161 N34160 N34161 10
D34161 N34161 0 diode
R34162 N34161 N34162 10
D34162 N34162 0 diode
R34163 N34162 N34163 10
D34163 N34163 0 diode
R34164 N34163 N34164 10
D34164 N34164 0 diode
R34165 N34164 N34165 10
D34165 N34165 0 diode
R34166 N34165 N34166 10
D34166 N34166 0 diode
R34167 N34166 N34167 10
D34167 N34167 0 diode
R34168 N34167 N34168 10
D34168 N34168 0 diode
R34169 N34168 N34169 10
D34169 N34169 0 diode
R34170 N34169 N34170 10
D34170 N34170 0 diode
R34171 N34170 N34171 10
D34171 N34171 0 diode
R34172 N34171 N34172 10
D34172 N34172 0 diode
R34173 N34172 N34173 10
D34173 N34173 0 diode
R34174 N34173 N34174 10
D34174 N34174 0 diode
R34175 N34174 N34175 10
D34175 N34175 0 diode
R34176 N34175 N34176 10
D34176 N34176 0 diode
R34177 N34176 N34177 10
D34177 N34177 0 diode
R34178 N34177 N34178 10
D34178 N34178 0 diode
R34179 N34178 N34179 10
D34179 N34179 0 diode
R34180 N34179 N34180 10
D34180 N34180 0 diode
R34181 N34180 N34181 10
D34181 N34181 0 diode
R34182 N34181 N34182 10
D34182 N34182 0 diode
R34183 N34182 N34183 10
D34183 N34183 0 diode
R34184 N34183 N34184 10
D34184 N34184 0 diode
R34185 N34184 N34185 10
D34185 N34185 0 diode
R34186 N34185 N34186 10
D34186 N34186 0 diode
R34187 N34186 N34187 10
D34187 N34187 0 diode
R34188 N34187 N34188 10
D34188 N34188 0 diode
R34189 N34188 N34189 10
D34189 N34189 0 diode
R34190 N34189 N34190 10
D34190 N34190 0 diode
R34191 N34190 N34191 10
D34191 N34191 0 diode
R34192 N34191 N34192 10
D34192 N34192 0 diode
R34193 N34192 N34193 10
D34193 N34193 0 diode
R34194 N34193 N34194 10
D34194 N34194 0 diode
R34195 N34194 N34195 10
D34195 N34195 0 diode
R34196 N34195 N34196 10
D34196 N34196 0 diode
R34197 N34196 N34197 10
D34197 N34197 0 diode
R34198 N34197 N34198 10
D34198 N34198 0 diode
R34199 N34198 N34199 10
D34199 N34199 0 diode
R34200 N34199 N34200 10
D34200 N34200 0 diode
R34201 N34200 N34201 10
D34201 N34201 0 diode
R34202 N34201 N34202 10
D34202 N34202 0 diode
R34203 N34202 N34203 10
D34203 N34203 0 diode
R34204 N34203 N34204 10
D34204 N34204 0 diode
R34205 N34204 N34205 10
D34205 N34205 0 diode
R34206 N34205 N34206 10
D34206 N34206 0 diode
R34207 N34206 N34207 10
D34207 N34207 0 diode
R34208 N34207 N34208 10
D34208 N34208 0 diode
R34209 N34208 N34209 10
D34209 N34209 0 diode
R34210 N34209 N34210 10
D34210 N34210 0 diode
R34211 N34210 N34211 10
D34211 N34211 0 diode
R34212 N34211 N34212 10
D34212 N34212 0 diode
R34213 N34212 N34213 10
D34213 N34213 0 diode
R34214 N34213 N34214 10
D34214 N34214 0 diode
R34215 N34214 N34215 10
D34215 N34215 0 diode
R34216 N34215 N34216 10
D34216 N34216 0 diode
R34217 N34216 N34217 10
D34217 N34217 0 diode
R34218 N34217 N34218 10
D34218 N34218 0 diode
R34219 N34218 N34219 10
D34219 N34219 0 diode
R34220 N34219 N34220 10
D34220 N34220 0 diode
R34221 N34220 N34221 10
D34221 N34221 0 diode
R34222 N34221 N34222 10
D34222 N34222 0 diode
R34223 N34222 N34223 10
D34223 N34223 0 diode
R34224 N34223 N34224 10
D34224 N34224 0 diode
R34225 N34224 N34225 10
D34225 N34225 0 diode
R34226 N34225 N34226 10
D34226 N34226 0 diode
R34227 N34226 N34227 10
D34227 N34227 0 diode
R34228 N34227 N34228 10
D34228 N34228 0 diode
R34229 N34228 N34229 10
D34229 N34229 0 diode
R34230 N34229 N34230 10
D34230 N34230 0 diode
R34231 N34230 N34231 10
D34231 N34231 0 diode
R34232 N34231 N34232 10
D34232 N34232 0 diode
R34233 N34232 N34233 10
D34233 N34233 0 diode
R34234 N34233 N34234 10
D34234 N34234 0 diode
R34235 N34234 N34235 10
D34235 N34235 0 diode
R34236 N34235 N34236 10
D34236 N34236 0 diode
R34237 N34236 N34237 10
D34237 N34237 0 diode
R34238 N34237 N34238 10
D34238 N34238 0 diode
R34239 N34238 N34239 10
D34239 N34239 0 diode
R34240 N34239 N34240 10
D34240 N34240 0 diode
R34241 N34240 N34241 10
D34241 N34241 0 diode
R34242 N34241 N34242 10
D34242 N34242 0 diode
R34243 N34242 N34243 10
D34243 N34243 0 diode
R34244 N34243 N34244 10
D34244 N34244 0 diode
R34245 N34244 N34245 10
D34245 N34245 0 diode
R34246 N34245 N34246 10
D34246 N34246 0 diode
R34247 N34246 N34247 10
D34247 N34247 0 diode
R34248 N34247 N34248 10
D34248 N34248 0 diode
R34249 N34248 N34249 10
D34249 N34249 0 diode
R34250 N34249 N34250 10
D34250 N34250 0 diode
R34251 N34250 N34251 10
D34251 N34251 0 diode
R34252 N34251 N34252 10
D34252 N34252 0 diode
R34253 N34252 N34253 10
D34253 N34253 0 diode
R34254 N34253 N34254 10
D34254 N34254 0 diode
R34255 N34254 N34255 10
D34255 N34255 0 diode
R34256 N34255 N34256 10
D34256 N34256 0 diode
R34257 N34256 N34257 10
D34257 N34257 0 diode
R34258 N34257 N34258 10
D34258 N34258 0 diode
R34259 N34258 N34259 10
D34259 N34259 0 diode
R34260 N34259 N34260 10
D34260 N34260 0 diode
R34261 N34260 N34261 10
D34261 N34261 0 diode
R34262 N34261 N34262 10
D34262 N34262 0 diode
R34263 N34262 N34263 10
D34263 N34263 0 diode
R34264 N34263 N34264 10
D34264 N34264 0 diode
R34265 N34264 N34265 10
D34265 N34265 0 diode
R34266 N34265 N34266 10
D34266 N34266 0 diode
R34267 N34266 N34267 10
D34267 N34267 0 diode
R34268 N34267 N34268 10
D34268 N34268 0 diode
R34269 N34268 N34269 10
D34269 N34269 0 diode
R34270 N34269 N34270 10
D34270 N34270 0 diode
R34271 N34270 N34271 10
D34271 N34271 0 diode
R34272 N34271 N34272 10
D34272 N34272 0 diode
R34273 N34272 N34273 10
D34273 N34273 0 diode
R34274 N34273 N34274 10
D34274 N34274 0 diode
R34275 N34274 N34275 10
D34275 N34275 0 diode
R34276 N34275 N34276 10
D34276 N34276 0 diode
R34277 N34276 N34277 10
D34277 N34277 0 diode
R34278 N34277 N34278 10
D34278 N34278 0 diode
R34279 N34278 N34279 10
D34279 N34279 0 diode
R34280 N34279 N34280 10
D34280 N34280 0 diode
R34281 N34280 N34281 10
D34281 N34281 0 diode
R34282 N34281 N34282 10
D34282 N34282 0 diode
R34283 N34282 N34283 10
D34283 N34283 0 diode
R34284 N34283 N34284 10
D34284 N34284 0 diode
R34285 N34284 N34285 10
D34285 N34285 0 diode
R34286 N34285 N34286 10
D34286 N34286 0 diode
R34287 N34286 N34287 10
D34287 N34287 0 diode
R34288 N34287 N34288 10
D34288 N34288 0 diode
R34289 N34288 N34289 10
D34289 N34289 0 diode
R34290 N34289 N34290 10
D34290 N34290 0 diode
R34291 N34290 N34291 10
D34291 N34291 0 diode
R34292 N34291 N34292 10
D34292 N34292 0 diode
R34293 N34292 N34293 10
D34293 N34293 0 diode
R34294 N34293 N34294 10
D34294 N34294 0 diode
R34295 N34294 N34295 10
D34295 N34295 0 diode
R34296 N34295 N34296 10
D34296 N34296 0 diode
R34297 N34296 N34297 10
D34297 N34297 0 diode
R34298 N34297 N34298 10
D34298 N34298 0 diode
R34299 N34298 N34299 10
D34299 N34299 0 diode
R34300 N34299 N34300 10
D34300 N34300 0 diode
R34301 N34300 N34301 10
D34301 N34301 0 diode
R34302 N34301 N34302 10
D34302 N34302 0 diode
R34303 N34302 N34303 10
D34303 N34303 0 diode
R34304 N34303 N34304 10
D34304 N34304 0 diode
R34305 N34304 N34305 10
D34305 N34305 0 diode
R34306 N34305 N34306 10
D34306 N34306 0 diode
R34307 N34306 N34307 10
D34307 N34307 0 diode
R34308 N34307 N34308 10
D34308 N34308 0 diode
R34309 N34308 N34309 10
D34309 N34309 0 diode
R34310 N34309 N34310 10
D34310 N34310 0 diode
R34311 N34310 N34311 10
D34311 N34311 0 diode
R34312 N34311 N34312 10
D34312 N34312 0 diode
R34313 N34312 N34313 10
D34313 N34313 0 diode
R34314 N34313 N34314 10
D34314 N34314 0 diode
R34315 N34314 N34315 10
D34315 N34315 0 diode
R34316 N34315 N34316 10
D34316 N34316 0 diode
R34317 N34316 N34317 10
D34317 N34317 0 diode
R34318 N34317 N34318 10
D34318 N34318 0 diode
R34319 N34318 N34319 10
D34319 N34319 0 diode
R34320 N34319 N34320 10
D34320 N34320 0 diode
R34321 N34320 N34321 10
D34321 N34321 0 diode
R34322 N34321 N34322 10
D34322 N34322 0 diode
R34323 N34322 N34323 10
D34323 N34323 0 diode
R34324 N34323 N34324 10
D34324 N34324 0 diode
R34325 N34324 N34325 10
D34325 N34325 0 diode
R34326 N34325 N34326 10
D34326 N34326 0 diode
R34327 N34326 N34327 10
D34327 N34327 0 diode
R34328 N34327 N34328 10
D34328 N34328 0 diode
R34329 N34328 N34329 10
D34329 N34329 0 diode
R34330 N34329 N34330 10
D34330 N34330 0 diode
R34331 N34330 N34331 10
D34331 N34331 0 diode
R34332 N34331 N34332 10
D34332 N34332 0 diode
R34333 N34332 N34333 10
D34333 N34333 0 diode
R34334 N34333 N34334 10
D34334 N34334 0 diode
R34335 N34334 N34335 10
D34335 N34335 0 diode
R34336 N34335 N34336 10
D34336 N34336 0 diode
R34337 N34336 N34337 10
D34337 N34337 0 diode
R34338 N34337 N34338 10
D34338 N34338 0 diode
R34339 N34338 N34339 10
D34339 N34339 0 diode
R34340 N34339 N34340 10
D34340 N34340 0 diode
R34341 N34340 N34341 10
D34341 N34341 0 diode
R34342 N34341 N34342 10
D34342 N34342 0 diode
R34343 N34342 N34343 10
D34343 N34343 0 diode
R34344 N34343 N34344 10
D34344 N34344 0 diode
R34345 N34344 N34345 10
D34345 N34345 0 diode
R34346 N34345 N34346 10
D34346 N34346 0 diode
R34347 N34346 N34347 10
D34347 N34347 0 diode
R34348 N34347 N34348 10
D34348 N34348 0 diode
R34349 N34348 N34349 10
D34349 N34349 0 diode
R34350 N34349 N34350 10
D34350 N34350 0 diode
R34351 N34350 N34351 10
D34351 N34351 0 diode
R34352 N34351 N34352 10
D34352 N34352 0 diode
R34353 N34352 N34353 10
D34353 N34353 0 diode
R34354 N34353 N34354 10
D34354 N34354 0 diode
R34355 N34354 N34355 10
D34355 N34355 0 diode
R34356 N34355 N34356 10
D34356 N34356 0 diode
R34357 N34356 N34357 10
D34357 N34357 0 diode
R34358 N34357 N34358 10
D34358 N34358 0 diode
R34359 N34358 N34359 10
D34359 N34359 0 diode
R34360 N34359 N34360 10
D34360 N34360 0 diode
R34361 N34360 N34361 10
D34361 N34361 0 diode
R34362 N34361 N34362 10
D34362 N34362 0 diode
R34363 N34362 N34363 10
D34363 N34363 0 diode
R34364 N34363 N34364 10
D34364 N34364 0 diode
R34365 N34364 N34365 10
D34365 N34365 0 diode
R34366 N34365 N34366 10
D34366 N34366 0 diode
R34367 N34366 N34367 10
D34367 N34367 0 diode
R34368 N34367 N34368 10
D34368 N34368 0 diode
R34369 N34368 N34369 10
D34369 N34369 0 diode
R34370 N34369 N34370 10
D34370 N34370 0 diode
R34371 N34370 N34371 10
D34371 N34371 0 diode
R34372 N34371 N34372 10
D34372 N34372 0 diode
R34373 N34372 N34373 10
D34373 N34373 0 diode
R34374 N34373 N34374 10
D34374 N34374 0 diode
R34375 N34374 N34375 10
D34375 N34375 0 diode
R34376 N34375 N34376 10
D34376 N34376 0 diode
R34377 N34376 N34377 10
D34377 N34377 0 diode
R34378 N34377 N34378 10
D34378 N34378 0 diode
R34379 N34378 N34379 10
D34379 N34379 0 diode
R34380 N34379 N34380 10
D34380 N34380 0 diode
R34381 N34380 N34381 10
D34381 N34381 0 diode
R34382 N34381 N34382 10
D34382 N34382 0 diode
R34383 N34382 N34383 10
D34383 N34383 0 diode
R34384 N34383 N34384 10
D34384 N34384 0 diode
R34385 N34384 N34385 10
D34385 N34385 0 diode
R34386 N34385 N34386 10
D34386 N34386 0 diode
R34387 N34386 N34387 10
D34387 N34387 0 diode
R34388 N34387 N34388 10
D34388 N34388 0 diode
R34389 N34388 N34389 10
D34389 N34389 0 diode
R34390 N34389 N34390 10
D34390 N34390 0 diode
R34391 N34390 N34391 10
D34391 N34391 0 diode
R34392 N34391 N34392 10
D34392 N34392 0 diode
R34393 N34392 N34393 10
D34393 N34393 0 diode
R34394 N34393 N34394 10
D34394 N34394 0 diode
R34395 N34394 N34395 10
D34395 N34395 0 diode
R34396 N34395 N34396 10
D34396 N34396 0 diode
R34397 N34396 N34397 10
D34397 N34397 0 diode
R34398 N34397 N34398 10
D34398 N34398 0 diode
R34399 N34398 N34399 10
D34399 N34399 0 diode
R34400 N34399 N34400 10
D34400 N34400 0 diode
R34401 N34400 N34401 10
D34401 N34401 0 diode
R34402 N34401 N34402 10
D34402 N34402 0 diode
R34403 N34402 N34403 10
D34403 N34403 0 diode
R34404 N34403 N34404 10
D34404 N34404 0 diode
R34405 N34404 N34405 10
D34405 N34405 0 diode
R34406 N34405 N34406 10
D34406 N34406 0 diode
R34407 N34406 N34407 10
D34407 N34407 0 diode
R34408 N34407 N34408 10
D34408 N34408 0 diode
R34409 N34408 N34409 10
D34409 N34409 0 diode
R34410 N34409 N34410 10
D34410 N34410 0 diode
R34411 N34410 N34411 10
D34411 N34411 0 diode
R34412 N34411 N34412 10
D34412 N34412 0 diode
R34413 N34412 N34413 10
D34413 N34413 0 diode
R34414 N34413 N34414 10
D34414 N34414 0 diode
R34415 N34414 N34415 10
D34415 N34415 0 diode
R34416 N34415 N34416 10
D34416 N34416 0 diode
R34417 N34416 N34417 10
D34417 N34417 0 diode
R34418 N34417 N34418 10
D34418 N34418 0 diode
R34419 N34418 N34419 10
D34419 N34419 0 diode
R34420 N34419 N34420 10
D34420 N34420 0 diode
R34421 N34420 N34421 10
D34421 N34421 0 diode
R34422 N34421 N34422 10
D34422 N34422 0 diode
R34423 N34422 N34423 10
D34423 N34423 0 diode
R34424 N34423 N34424 10
D34424 N34424 0 diode
R34425 N34424 N34425 10
D34425 N34425 0 diode
R34426 N34425 N34426 10
D34426 N34426 0 diode
R34427 N34426 N34427 10
D34427 N34427 0 diode
R34428 N34427 N34428 10
D34428 N34428 0 diode
R34429 N34428 N34429 10
D34429 N34429 0 diode
R34430 N34429 N34430 10
D34430 N34430 0 diode
R34431 N34430 N34431 10
D34431 N34431 0 diode
R34432 N34431 N34432 10
D34432 N34432 0 diode
R34433 N34432 N34433 10
D34433 N34433 0 diode
R34434 N34433 N34434 10
D34434 N34434 0 diode
R34435 N34434 N34435 10
D34435 N34435 0 diode
R34436 N34435 N34436 10
D34436 N34436 0 diode
R34437 N34436 N34437 10
D34437 N34437 0 diode
R34438 N34437 N34438 10
D34438 N34438 0 diode
R34439 N34438 N34439 10
D34439 N34439 0 diode
R34440 N34439 N34440 10
D34440 N34440 0 diode
R34441 N34440 N34441 10
D34441 N34441 0 diode
R34442 N34441 N34442 10
D34442 N34442 0 diode
R34443 N34442 N34443 10
D34443 N34443 0 diode
R34444 N34443 N34444 10
D34444 N34444 0 diode
R34445 N34444 N34445 10
D34445 N34445 0 diode
R34446 N34445 N34446 10
D34446 N34446 0 diode
R34447 N34446 N34447 10
D34447 N34447 0 diode
R34448 N34447 N34448 10
D34448 N34448 0 diode
R34449 N34448 N34449 10
D34449 N34449 0 diode
R34450 N34449 N34450 10
D34450 N34450 0 diode
R34451 N34450 N34451 10
D34451 N34451 0 diode
R34452 N34451 N34452 10
D34452 N34452 0 diode
R34453 N34452 N34453 10
D34453 N34453 0 diode
R34454 N34453 N34454 10
D34454 N34454 0 diode
R34455 N34454 N34455 10
D34455 N34455 0 diode
R34456 N34455 N34456 10
D34456 N34456 0 diode
R34457 N34456 N34457 10
D34457 N34457 0 diode
R34458 N34457 N34458 10
D34458 N34458 0 diode
R34459 N34458 N34459 10
D34459 N34459 0 diode
R34460 N34459 N34460 10
D34460 N34460 0 diode
R34461 N34460 N34461 10
D34461 N34461 0 diode
R34462 N34461 N34462 10
D34462 N34462 0 diode
R34463 N34462 N34463 10
D34463 N34463 0 diode
R34464 N34463 N34464 10
D34464 N34464 0 diode
R34465 N34464 N34465 10
D34465 N34465 0 diode
R34466 N34465 N34466 10
D34466 N34466 0 diode
R34467 N34466 N34467 10
D34467 N34467 0 diode
R34468 N34467 N34468 10
D34468 N34468 0 diode
R34469 N34468 N34469 10
D34469 N34469 0 diode
R34470 N34469 N34470 10
D34470 N34470 0 diode
R34471 N34470 N34471 10
D34471 N34471 0 diode
R34472 N34471 N34472 10
D34472 N34472 0 diode
R34473 N34472 N34473 10
D34473 N34473 0 diode
R34474 N34473 N34474 10
D34474 N34474 0 diode
R34475 N34474 N34475 10
D34475 N34475 0 diode
R34476 N34475 N34476 10
D34476 N34476 0 diode
R34477 N34476 N34477 10
D34477 N34477 0 diode
R34478 N34477 N34478 10
D34478 N34478 0 diode
R34479 N34478 N34479 10
D34479 N34479 0 diode
R34480 N34479 N34480 10
D34480 N34480 0 diode
R34481 N34480 N34481 10
D34481 N34481 0 diode
R34482 N34481 N34482 10
D34482 N34482 0 diode
R34483 N34482 N34483 10
D34483 N34483 0 diode
R34484 N34483 N34484 10
D34484 N34484 0 diode
R34485 N34484 N34485 10
D34485 N34485 0 diode
R34486 N34485 N34486 10
D34486 N34486 0 diode
R34487 N34486 N34487 10
D34487 N34487 0 diode
R34488 N34487 N34488 10
D34488 N34488 0 diode
R34489 N34488 N34489 10
D34489 N34489 0 diode
R34490 N34489 N34490 10
D34490 N34490 0 diode
R34491 N34490 N34491 10
D34491 N34491 0 diode
R34492 N34491 N34492 10
D34492 N34492 0 diode
R34493 N34492 N34493 10
D34493 N34493 0 diode
R34494 N34493 N34494 10
D34494 N34494 0 diode
R34495 N34494 N34495 10
D34495 N34495 0 diode
R34496 N34495 N34496 10
D34496 N34496 0 diode
R34497 N34496 N34497 10
D34497 N34497 0 diode
R34498 N34497 N34498 10
D34498 N34498 0 diode
R34499 N34498 N34499 10
D34499 N34499 0 diode
R34500 N34499 N34500 10
D34500 N34500 0 diode
R34501 N34500 N34501 10
D34501 N34501 0 diode
R34502 N34501 N34502 10
D34502 N34502 0 diode
R34503 N34502 N34503 10
D34503 N34503 0 diode
R34504 N34503 N34504 10
D34504 N34504 0 diode
R34505 N34504 N34505 10
D34505 N34505 0 diode
R34506 N34505 N34506 10
D34506 N34506 0 diode
R34507 N34506 N34507 10
D34507 N34507 0 diode
R34508 N34507 N34508 10
D34508 N34508 0 diode
R34509 N34508 N34509 10
D34509 N34509 0 diode
R34510 N34509 N34510 10
D34510 N34510 0 diode
R34511 N34510 N34511 10
D34511 N34511 0 diode
R34512 N34511 N34512 10
D34512 N34512 0 diode
R34513 N34512 N34513 10
D34513 N34513 0 diode
R34514 N34513 N34514 10
D34514 N34514 0 diode
R34515 N34514 N34515 10
D34515 N34515 0 diode
R34516 N34515 N34516 10
D34516 N34516 0 diode
R34517 N34516 N34517 10
D34517 N34517 0 diode
R34518 N34517 N34518 10
D34518 N34518 0 diode
R34519 N34518 N34519 10
D34519 N34519 0 diode
R34520 N34519 N34520 10
D34520 N34520 0 diode
R34521 N34520 N34521 10
D34521 N34521 0 diode
R34522 N34521 N34522 10
D34522 N34522 0 diode
R34523 N34522 N34523 10
D34523 N34523 0 diode
R34524 N34523 N34524 10
D34524 N34524 0 diode
R34525 N34524 N34525 10
D34525 N34525 0 diode
R34526 N34525 N34526 10
D34526 N34526 0 diode
R34527 N34526 N34527 10
D34527 N34527 0 diode
R34528 N34527 N34528 10
D34528 N34528 0 diode
R34529 N34528 N34529 10
D34529 N34529 0 diode
R34530 N34529 N34530 10
D34530 N34530 0 diode
R34531 N34530 N34531 10
D34531 N34531 0 diode
R34532 N34531 N34532 10
D34532 N34532 0 diode
R34533 N34532 N34533 10
D34533 N34533 0 diode
R34534 N34533 N34534 10
D34534 N34534 0 diode
R34535 N34534 N34535 10
D34535 N34535 0 diode
R34536 N34535 N34536 10
D34536 N34536 0 diode
R34537 N34536 N34537 10
D34537 N34537 0 diode
R34538 N34537 N34538 10
D34538 N34538 0 diode
R34539 N34538 N34539 10
D34539 N34539 0 diode
R34540 N34539 N34540 10
D34540 N34540 0 diode
R34541 N34540 N34541 10
D34541 N34541 0 diode
R34542 N34541 N34542 10
D34542 N34542 0 diode
R34543 N34542 N34543 10
D34543 N34543 0 diode
R34544 N34543 N34544 10
D34544 N34544 0 diode
R34545 N34544 N34545 10
D34545 N34545 0 diode
R34546 N34545 N34546 10
D34546 N34546 0 diode
R34547 N34546 N34547 10
D34547 N34547 0 diode
R34548 N34547 N34548 10
D34548 N34548 0 diode
R34549 N34548 N34549 10
D34549 N34549 0 diode
R34550 N34549 N34550 10
D34550 N34550 0 diode
R34551 N34550 N34551 10
D34551 N34551 0 diode
R34552 N34551 N34552 10
D34552 N34552 0 diode
R34553 N34552 N34553 10
D34553 N34553 0 diode
R34554 N34553 N34554 10
D34554 N34554 0 diode
R34555 N34554 N34555 10
D34555 N34555 0 diode
R34556 N34555 N34556 10
D34556 N34556 0 diode
R34557 N34556 N34557 10
D34557 N34557 0 diode
R34558 N34557 N34558 10
D34558 N34558 0 diode
R34559 N34558 N34559 10
D34559 N34559 0 diode
R34560 N34559 N34560 10
D34560 N34560 0 diode
R34561 N34560 N34561 10
D34561 N34561 0 diode
R34562 N34561 N34562 10
D34562 N34562 0 diode
R34563 N34562 N34563 10
D34563 N34563 0 diode
R34564 N34563 N34564 10
D34564 N34564 0 diode
R34565 N34564 N34565 10
D34565 N34565 0 diode
R34566 N34565 N34566 10
D34566 N34566 0 diode
R34567 N34566 N34567 10
D34567 N34567 0 diode
R34568 N34567 N34568 10
D34568 N34568 0 diode
R34569 N34568 N34569 10
D34569 N34569 0 diode
R34570 N34569 N34570 10
D34570 N34570 0 diode
R34571 N34570 N34571 10
D34571 N34571 0 diode
R34572 N34571 N34572 10
D34572 N34572 0 diode
R34573 N34572 N34573 10
D34573 N34573 0 diode
R34574 N34573 N34574 10
D34574 N34574 0 diode
R34575 N34574 N34575 10
D34575 N34575 0 diode
R34576 N34575 N34576 10
D34576 N34576 0 diode
R34577 N34576 N34577 10
D34577 N34577 0 diode
R34578 N34577 N34578 10
D34578 N34578 0 diode
R34579 N34578 N34579 10
D34579 N34579 0 diode
R34580 N34579 N34580 10
D34580 N34580 0 diode
R34581 N34580 N34581 10
D34581 N34581 0 diode
R34582 N34581 N34582 10
D34582 N34582 0 diode
R34583 N34582 N34583 10
D34583 N34583 0 diode
R34584 N34583 N34584 10
D34584 N34584 0 diode
R34585 N34584 N34585 10
D34585 N34585 0 diode
R34586 N34585 N34586 10
D34586 N34586 0 diode
R34587 N34586 N34587 10
D34587 N34587 0 diode
R34588 N34587 N34588 10
D34588 N34588 0 diode
R34589 N34588 N34589 10
D34589 N34589 0 diode
R34590 N34589 N34590 10
D34590 N34590 0 diode
R34591 N34590 N34591 10
D34591 N34591 0 diode
R34592 N34591 N34592 10
D34592 N34592 0 diode
R34593 N34592 N34593 10
D34593 N34593 0 diode
R34594 N34593 N34594 10
D34594 N34594 0 diode
R34595 N34594 N34595 10
D34595 N34595 0 diode
R34596 N34595 N34596 10
D34596 N34596 0 diode
R34597 N34596 N34597 10
D34597 N34597 0 diode
R34598 N34597 N34598 10
D34598 N34598 0 diode
R34599 N34598 N34599 10
D34599 N34599 0 diode
R34600 N34599 N34600 10
D34600 N34600 0 diode
R34601 N34600 N34601 10
D34601 N34601 0 diode
R34602 N34601 N34602 10
D34602 N34602 0 diode
R34603 N34602 N34603 10
D34603 N34603 0 diode
R34604 N34603 N34604 10
D34604 N34604 0 diode
R34605 N34604 N34605 10
D34605 N34605 0 diode
R34606 N34605 N34606 10
D34606 N34606 0 diode
R34607 N34606 N34607 10
D34607 N34607 0 diode
R34608 N34607 N34608 10
D34608 N34608 0 diode
R34609 N34608 N34609 10
D34609 N34609 0 diode
R34610 N34609 N34610 10
D34610 N34610 0 diode
R34611 N34610 N34611 10
D34611 N34611 0 diode
R34612 N34611 N34612 10
D34612 N34612 0 diode
R34613 N34612 N34613 10
D34613 N34613 0 diode
R34614 N34613 N34614 10
D34614 N34614 0 diode
R34615 N34614 N34615 10
D34615 N34615 0 diode
R34616 N34615 N34616 10
D34616 N34616 0 diode
R34617 N34616 N34617 10
D34617 N34617 0 diode
R34618 N34617 N34618 10
D34618 N34618 0 diode
R34619 N34618 N34619 10
D34619 N34619 0 diode
R34620 N34619 N34620 10
D34620 N34620 0 diode
R34621 N34620 N34621 10
D34621 N34621 0 diode
R34622 N34621 N34622 10
D34622 N34622 0 diode
R34623 N34622 N34623 10
D34623 N34623 0 diode
R34624 N34623 N34624 10
D34624 N34624 0 diode
R34625 N34624 N34625 10
D34625 N34625 0 diode
R34626 N34625 N34626 10
D34626 N34626 0 diode
R34627 N34626 N34627 10
D34627 N34627 0 diode
R34628 N34627 N34628 10
D34628 N34628 0 diode
R34629 N34628 N34629 10
D34629 N34629 0 diode
R34630 N34629 N34630 10
D34630 N34630 0 diode
R34631 N34630 N34631 10
D34631 N34631 0 diode
R34632 N34631 N34632 10
D34632 N34632 0 diode
R34633 N34632 N34633 10
D34633 N34633 0 diode
R34634 N34633 N34634 10
D34634 N34634 0 diode
R34635 N34634 N34635 10
D34635 N34635 0 diode
R34636 N34635 N34636 10
D34636 N34636 0 diode
R34637 N34636 N34637 10
D34637 N34637 0 diode
R34638 N34637 N34638 10
D34638 N34638 0 diode
R34639 N34638 N34639 10
D34639 N34639 0 diode
R34640 N34639 N34640 10
D34640 N34640 0 diode
R34641 N34640 N34641 10
D34641 N34641 0 diode
R34642 N34641 N34642 10
D34642 N34642 0 diode
R34643 N34642 N34643 10
D34643 N34643 0 diode
R34644 N34643 N34644 10
D34644 N34644 0 diode
R34645 N34644 N34645 10
D34645 N34645 0 diode
R34646 N34645 N34646 10
D34646 N34646 0 diode
R34647 N34646 N34647 10
D34647 N34647 0 diode
R34648 N34647 N34648 10
D34648 N34648 0 diode
R34649 N34648 N34649 10
D34649 N34649 0 diode
R34650 N34649 N34650 10
D34650 N34650 0 diode
R34651 N34650 N34651 10
D34651 N34651 0 diode
R34652 N34651 N34652 10
D34652 N34652 0 diode
R34653 N34652 N34653 10
D34653 N34653 0 diode
R34654 N34653 N34654 10
D34654 N34654 0 diode
R34655 N34654 N34655 10
D34655 N34655 0 diode
R34656 N34655 N34656 10
D34656 N34656 0 diode
R34657 N34656 N34657 10
D34657 N34657 0 diode
R34658 N34657 N34658 10
D34658 N34658 0 diode
R34659 N34658 N34659 10
D34659 N34659 0 diode
R34660 N34659 N34660 10
D34660 N34660 0 diode
R34661 N34660 N34661 10
D34661 N34661 0 diode
R34662 N34661 N34662 10
D34662 N34662 0 diode
R34663 N34662 N34663 10
D34663 N34663 0 diode
R34664 N34663 N34664 10
D34664 N34664 0 diode
R34665 N34664 N34665 10
D34665 N34665 0 diode
R34666 N34665 N34666 10
D34666 N34666 0 diode
R34667 N34666 N34667 10
D34667 N34667 0 diode
R34668 N34667 N34668 10
D34668 N34668 0 diode
R34669 N34668 N34669 10
D34669 N34669 0 diode
R34670 N34669 N34670 10
D34670 N34670 0 diode
R34671 N34670 N34671 10
D34671 N34671 0 diode
R34672 N34671 N34672 10
D34672 N34672 0 diode
R34673 N34672 N34673 10
D34673 N34673 0 diode
R34674 N34673 N34674 10
D34674 N34674 0 diode
R34675 N34674 N34675 10
D34675 N34675 0 diode
R34676 N34675 N34676 10
D34676 N34676 0 diode
R34677 N34676 N34677 10
D34677 N34677 0 diode
R34678 N34677 N34678 10
D34678 N34678 0 diode
R34679 N34678 N34679 10
D34679 N34679 0 diode
R34680 N34679 N34680 10
D34680 N34680 0 diode
R34681 N34680 N34681 10
D34681 N34681 0 diode
R34682 N34681 N34682 10
D34682 N34682 0 diode
R34683 N34682 N34683 10
D34683 N34683 0 diode
R34684 N34683 N34684 10
D34684 N34684 0 diode
R34685 N34684 N34685 10
D34685 N34685 0 diode
R34686 N34685 N34686 10
D34686 N34686 0 diode
R34687 N34686 N34687 10
D34687 N34687 0 diode
R34688 N34687 N34688 10
D34688 N34688 0 diode
R34689 N34688 N34689 10
D34689 N34689 0 diode
R34690 N34689 N34690 10
D34690 N34690 0 diode
R34691 N34690 N34691 10
D34691 N34691 0 diode
R34692 N34691 N34692 10
D34692 N34692 0 diode
R34693 N34692 N34693 10
D34693 N34693 0 diode
R34694 N34693 N34694 10
D34694 N34694 0 diode
R34695 N34694 N34695 10
D34695 N34695 0 diode
R34696 N34695 N34696 10
D34696 N34696 0 diode
R34697 N34696 N34697 10
D34697 N34697 0 diode
R34698 N34697 N34698 10
D34698 N34698 0 diode
R34699 N34698 N34699 10
D34699 N34699 0 diode
R34700 N34699 N34700 10
D34700 N34700 0 diode
R34701 N34700 N34701 10
D34701 N34701 0 diode
R34702 N34701 N34702 10
D34702 N34702 0 diode
R34703 N34702 N34703 10
D34703 N34703 0 diode
R34704 N34703 N34704 10
D34704 N34704 0 diode
R34705 N34704 N34705 10
D34705 N34705 0 diode
R34706 N34705 N34706 10
D34706 N34706 0 diode
R34707 N34706 N34707 10
D34707 N34707 0 diode
R34708 N34707 N34708 10
D34708 N34708 0 diode
R34709 N34708 N34709 10
D34709 N34709 0 diode
R34710 N34709 N34710 10
D34710 N34710 0 diode
R34711 N34710 N34711 10
D34711 N34711 0 diode
R34712 N34711 N34712 10
D34712 N34712 0 diode
R34713 N34712 N34713 10
D34713 N34713 0 diode
R34714 N34713 N34714 10
D34714 N34714 0 diode
R34715 N34714 N34715 10
D34715 N34715 0 diode
R34716 N34715 N34716 10
D34716 N34716 0 diode
R34717 N34716 N34717 10
D34717 N34717 0 diode
R34718 N34717 N34718 10
D34718 N34718 0 diode
R34719 N34718 N34719 10
D34719 N34719 0 diode
R34720 N34719 N34720 10
D34720 N34720 0 diode
R34721 N34720 N34721 10
D34721 N34721 0 diode
R34722 N34721 N34722 10
D34722 N34722 0 diode
R34723 N34722 N34723 10
D34723 N34723 0 diode
R34724 N34723 N34724 10
D34724 N34724 0 diode
R34725 N34724 N34725 10
D34725 N34725 0 diode
R34726 N34725 N34726 10
D34726 N34726 0 diode
R34727 N34726 N34727 10
D34727 N34727 0 diode
R34728 N34727 N34728 10
D34728 N34728 0 diode
R34729 N34728 N34729 10
D34729 N34729 0 diode
R34730 N34729 N34730 10
D34730 N34730 0 diode
R34731 N34730 N34731 10
D34731 N34731 0 diode
R34732 N34731 N34732 10
D34732 N34732 0 diode
R34733 N34732 N34733 10
D34733 N34733 0 diode
R34734 N34733 N34734 10
D34734 N34734 0 diode
R34735 N34734 N34735 10
D34735 N34735 0 diode
R34736 N34735 N34736 10
D34736 N34736 0 diode
R34737 N34736 N34737 10
D34737 N34737 0 diode
R34738 N34737 N34738 10
D34738 N34738 0 diode
R34739 N34738 N34739 10
D34739 N34739 0 diode
R34740 N34739 N34740 10
D34740 N34740 0 diode
R34741 N34740 N34741 10
D34741 N34741 0 diode
R34742 N34741 N34742 10
D34742 N34742 0 diode
R34743 N34742 N34743 10
D34743 N34743 0 diode
R34744 N34743 N34744 10
D34744 N34744 0 diode
R34745 N34744 N34745 10
D34745 N34745 0 diode
R34746 N34745 N34746 10
D34746 N34746 0 diode
R34747 N34746 N34747 10
D34747 N34747 0 diode
R34748 N34747 N34748 10
D34748 N34748 0 diode
R34749 N34748 N34749 10
D34749 N34749 0 diode
R34750 N34749 N34750 10
D34750 N34750 0 diode
R34751 N34750 N34751 10
D34751 N34751 0 diode
R34752 N34751 N34752 10
D34752 N34752 0 diode
R34753 N34752 N34753 10
D34753 N34753 0 diode
R34754 N34753 N34754 10
D34754 N34754 0 diode
R34755 N34754 N34755 10
D34755 N34755 0 diode
R34756 N34755 N34756 10
D34756 N34756 0 diode
R34757 N34756 N34757 10
D34757 N34757 0 diode
R34758 N34757 N34758 10
D34758 N34758 0 diode
R34759 N34758 N34759 10
D34759 N34759 0 diode
R34760 N34759 N34760 10
D34760 N34760 0 diode
R34761 N34760 N34761 10
D34761 N34761 0 diode
R34762 N34761 N34762 10
D34762 N34762 0 diode
R34763 N34762 N34763 10
D34763 N34763 0 diode
R34764 N34763 N34764 10
D34764 N34764 0 diode
R34765 N34764 N34765 10
D34765 N34765 0 diode
R34766 N34765 N34766 10
D34766 N34766 0 diode
R34767 N34766 N34767 10
D34767 N34767 0 diode
R34768 N34767 N34768 10
D34768 N34768 0 diode
R34769 N34768 N34769 10
D34769 N34769 0 diode
R34770 N34769 N34770 10
D34770 N34770 0 diode
R34771 N34770 N34771 10
D34771 N34771 0 diode
R34772 N34771 N34772 10
D34772 N34772 0 diode
R34773 N34772 N34773 10
D34773 N34773 0 diode
R34774 N34773 N34774 10
D34774 N34774 0 diode
R34775 N34774 N34775 10
D34775 N34775 0 diode
R34776 N34775 N34776 10
D34776 N34776 0 diode
R34777 N34776 N34777 10
D34777 N34777 0 diode
R34778 N34777 N34778 10
D34778 N34778 0 diode
R34779 N34778 N34779 10
D34779 N34779 0 diode
R34780 N34779 N34780 10
D34780 N34780 0 diode
R34781 N34780 N34781 10
D34781 N34781 0 diode
R34782 N34781 N34782 10
D34782 N34782 0 diode
R34783 N34782 N34783 10
D34783 N34783 0 diode
R34784 N34783 N34784 10
D34784 N34784 0 diode
R34785 N34784 N34785 10
D34785 N34785 0 diode
R34786 N34785 N34786 10
D34786 N34786 0 diode
R34787 N34786 N34787 10
D34787 N34787 0 diode
R34788 N34787 N34788 10
D34788 N34788 0 diode
R34789 N34788 N34789 10
D34789 N34789 0 diode
R34790 N34789 N34790 10
D34790 N34790 0 diode
R34791 N34790 N34791 10
D34791 N34791 0 diode
R34792 N34791 N34792 10
D34792 N34792 0 diode
R34793 N34792 N34793 10
D34793 N34793 0 diode
R34794 N34793 N34794 10
D34794 N34794 0 diode
R34795 N34794 N34795 10
D34795 N34795 0 diode
R34796 N34795 N34796 10
D34796 N34796 0 diode
R34797 N34796 N34797 10
D34797 N34797 0 diode
R34798 N34797 N34798 10
D34798 N34798 0 diode
R34799 N34798 N34799 10
D34799 N34799 0 diode
R34800 N34799 N34800 10
D34800 N34800 0 diode
R34801 N34800 N34801 10
D34801 N34801 0 diode
R34802 N34801 N34802 10
D34802 N34802 0 diode
R34803 N34802 N34803 10
D34803 N34803 0 diode
R34804 N34803 N34804 10
D34804 N34804 0 diode
R34805 N34804 N34805 10
D34805 N34805 0 diode
R34806 N34805 N34806 10
D34806 N34806 0 diode
R34807 N34806 N34807 10
D34807 N34807 0 diode
R34808 N34807 N34808 10
D34808 N34808 0 diode
R34809 N34808 N34809 10
D34809 N34809 0 diode
R34810 N34809 N34810 10
D34810 N34810 0 diode
R34811 N34810 N34811 10
D34811 N34811 0 diode
R34812 N34811 N34812 10
D34812 N34812 0 diode
R34813 N34812 N34813 10
D34813 N34813 0 diode
R34814 N34813 N34814 10
D34814 N34814 0 diode
R34815 N34814 N34815 10
D34815 N34815 0 diode
R34816 N34815 N34816 10
D34816 N34816 0 diode
R34817 N34816 N34817 10
D34817 N34817 0 diode
R34818 N34817 N34818 10
D34818 N34818 0 diode
R34819 N34818 N34819 10
D34819 N34819 0 diode
R34820 N34819 N34820 10
D34820 N34820 0 diode
R34821 N34820 N34821 10
D34821 N34821 0 diode
R34822 N34821 N34822 10
D34822 N34822 0 diode
R34823 N34822 N34823 10
D34823 N34823 0 diode
R34824 N34823 N34824 10
D34824 N34824 0 diode
R34825 N34824 N34825 10
D34825 N34825 0 diode
R34826 N34825 N34826 10
D34826 N34826 0 diode
R34827 N34826 N34827 10
D34827 N34827 0 diode
R34828 N34827 N34828 10
D34828 N34828 0 diode
R34829 N34828 N34829 10
D34829 N34829 0 diode
R34830 N34829 N34830 10
D34830 N34830 0 diode
R34831 N34830 N34831 10
D34831 N34831 0 diode
R34832 N34831 N34832 10
D34832 N34832 0 diode
R34833 N34832 N34833 10
D34833 N34833 0 diode
R34834 N34833 N34834 10
D34834 N34834 0 diode
R34835 N34834 N34835 10
D34835 N34835 0 diode
R34836 N34835 N34836 10
D34836 N34836 0 diode
R34837 N34836 N34837 10
D34837 N34837 0 diode
R34838 N34837 N34838 10
D34838 N34838 0 diode
R34839 N34838 N34839 10
D34839 N34839 0 diode
R34840 N34839 N34840 10
D34840 N34840 0 diode
R34841 N34840 N34841 10
D34841 N34841 0 diode
R34842 N34841 N34842 10
D34842 N34842 0 diode
R34843 N34842 N34843 10
D34843 N34843 0 diode
R34844 N34843 N34844 10
D34844 N34844 0 diode
R34845 N34844 N34845 10
D34845 N34845 0 diode
R34846 N34845 N34846 10
D34846 N34846 0 diode
R34847 N34846 N34847 10
D34847 N34847 0 diode
R34848 N34847 N34848 10
D34848 N34848 0 diode
R34849 N34848 N34849 10
D34849 N34849 0 diode
R34850 N34849 N34850 10
D34850 N34850 0 diode
R34851 N34850 N34851 10
D34851 N34851 0 diode
R34852 N34851 N34852 10
D34852 N34852 0 diode
R34853 N34852 N34853 10
D34853 N34853 0 diode
R34854 N34853 N34854 10
D34854 N34854 0 diode
R34855 N34854 N34855 10
D34855 N34855 0 diode
R34856 N34855 N34856 10
D34856 N34856 0 diode
R34857 N34856 N34857 10
D34857 N34857 0 diode
R34858 N34857 N34858 10
D34858 N34858 0 diode
R34859 N34858 N34859 10
D34859 N34859 0 diode
R34860 N34859 N34860 10
D34860 N34860 0 diode
R34861 N34860 N34861 10
D34861 N34861 0 diode
R34862 N34861 N34862 10
D34862 N34862 0 diode
R34863 N34862 N34863 10
D34863 N34863 0 diode
R34864 N34863 N34864 10
D34864 N34864 0 diode
R34865 N34864 N34865 10
D34865 N34865 0 diode
R34866 N34865 N34866 10
D34866 N34866 0 diode
R34867 N34866 N34867 10
D34867 N34867 0 diode
R34868 N34867 N34868 10
D34868 N34868 0 diode
R34869 N34868 N34869 10
D34869 N34869 0 diode
R34870 N34869 N34870 10
D34870 N34870 0 diode
R34871 N34870 N34871 10
D34871 N34871 0 diode
R34872 N34871 N34872 10
D34872 N34872 0 diode
R34873 N34872 N34873 10
D34873 N34873 0 diode
R34874 N34873 N34874 10
D34874 N34874 0 diode
R34875 N34874 N34875 10
D34875 N34875 0 diode
R34876 N34875 N34876 10
D34876 N34876 0 diode
R34877 N34876 N34877 10
D34877 N34877 0 diode
R34878 N34877 N34878 10
D34878 N34878 0 diode
R34879 N34878 N34879 10
D34879 N34879 0 diode
R34880 N34879 N34880 10
D34880 N34880 0 diode
R34881 N34880 N34881 10
D34881 N34881 0 diode
R34882 N34881 N34882 10
D34882 N34882 0 diode
R34883 N34882 N34883 10
D34883 N34883 0 diode
R34884 N34883 N34884 10
D34884 N34884 0 diode
R34885 N34884 N34885 10
D34885 N34885 0 diode
R34886 N34885 N34886 10
D34886 N34886 0 diode
R34887 N34886 N34887 10
D34887 N34887 0 diode
R34888 N34887 N34888 10
D34888 N34888 0 diode
R34889 N34888 N34889 10
D34889 N34889 0 diode
R34890 N34889 N34890 10
D34890 N34890 0 diode
R34891 N34890 N34891 10
D34891 N34891 0 diode
R34892 N34891 N34892 10
D34892 N34892 0 diode
R34893 N34892 N34893 10
D34893 N34893 0 diode
R34894 N34893 N34894 10
D34894 N34894 0 diode
R34895 N34894 N34895 10
D34895 N34895 0 diode
R34896 N34895 N34896 10
D34896 N34896 0 diode
R34897 N34896 N34897 10
D34897 N34897 0 diode
R34898 N34897 N34898 10
D34898 N34898 0 diode
R34899 N34898 N34899 10
D34899 N34899 0 diode
R34900 N34899 N34900 10
D34900 N34900 0 diode
R34901 N34900 N34901 10
D34901 N34901 0 diode
R34902 N34901 N34902 10
D34902 N34902 0 diode
R34903 N34902 N34903 10
D34903 N34903 0 diode
R34904 N34903 N34904 10
D34904 N34904 0 diode
R34905 N34904 N34905 10
D34905 N34905 0 diode
R34906 N34905 N34906 10
D34906 N34906 0 diode
R34907 N34906 N34907 10
D34907 N34907 0 diode
R34908 N34907 N34908 10
D34908 N34908 0 diode
R34909 N34908 N34909 10
D34909 N34909 0 diode
R34910 N34909 N34910 10
D34910 N34910 0 diode
R34911 N34910 N34911 10
D34911 N34911 0 diode
R34912 N34911 N34912 10
D34912 N34912 0 diode
R34913 N34912 N34913 10
D34913 N34913 0 diode
R34914 N34913 N34914 10
D34914 N34914 0 diode
R34915 N34914 N34915 10
D34915 N34915 0 diode
R34916 N34915 N34916 10
D34916 N34916 0 diode
R34917 N34916 N34917 10
D34917 N34917 0 diode
R34918 N34917 N34918 10
D34918 N34918 0 diode
R34919 N34918 N34919 10
D34919 N34919 0 diode
R34920 N34919 N34920 10
D34920 N34920 0 diode
R34921 N34920 N34921 10
D34921 N34921 0 diode
R34922 N34921 N34922 10
D34922 N34922 0 diode
R34923 N34922 N34923 10
D34923 N34923 0 diode
R34924 N34923 N34924 10
D34924 N34924 0 diode
R34925 N34924 N34925 10
D34925 N34925 0 diode
R34926 N34925 N34926 10
D34926 N34926 0 diode
R34927 N34926 N34927 10
D34927 N34927 0 diode
R34928 N34927 N34928 10
D34928 N34928 0 diode
R34929 N34928 N34929 10
D34929 N34929 0 diode
R34930 N34929 N34930 10
D34930 N34930 0 diode
R34931 N34930 N34931 10
D34931 N34931 0 diode
R34932 N34931 N34932 10
D34932 N34932 0 diode
R34933 N34932 N34933 10
D34933 N34933 0 diode
R34934 N34933 N34934 10
D34934 N34934 0 diode
R34935 N34934 N34935 10
D34935 N34935 0 diode
R34936 N34935 N34936 10
D34936 N34936 0 diode
R34937 N34936 N34937 10
D34937 N34937 0 diode
R34938 N34937 N34938 10
D34938 N34938 0 diode
R34939 N34938 N34939 10
D34939 N34939 0 diode
R34940 N34939 N34940 10
D34940 N34940 0 diode
R34941 N34940 N34941 10
D34941 N34941 0 diode
R34942 N34941 N34942 10
D34942 N34942 0 diode
R34943 N34942 N34943 10
D34943 N34943 0 diode
R34944 N34943 N34944 10
D34944 N34944 0 diode
R34945 N34944 N34945 10
D34945 N34945 0 diode
R34946 N34945 N34946 10
D34946 N34946 0 diode
R34947 N34946 N34947 10
D34947 N34947 0 diode
R34948 N34947 N34948 10
D34948 N34948 0 diode
R34949 N34948 N34949 10
D34949 N34949 0 diode
R34950 N34949 N34950 10
D34950 N34950 0 diode
R34951 N34950 N34951 10
D34951 N34951 0 diode
R34952 N34951 N34952 10
D34952 N34952 0 diode
R34953 N34952 N34953 10
D34953 N34953 0 diode
R34954 N34953 N34954 10
D34954 N34954 0 diode
R34955 N34954 N34955 10
D34955 N34955 0 diode
R34956 N34955 N34956 10
D34956 N34956 0 diode
R34957 N34956 N34957 10
D34957 N34957 0 diode
R34958 N34957 N34958 10
D34958 N34958 0 diode
R34959 N34958 N34959 10
D34959 N34959 0 diode
R34960 N34959 N34960 10
D34960 N34960 0 diode
R34961 N34960 N34961 10
D34961 N34961 0 diode
R34962 N34961 N34962 10
D34962 N34962 0 diode
R34963 N34962 N34963 10
D34963 N34963 0 diode
R34964 N34963 N34964 10
D34964 N34964 0 diode
R34965 N34964 N34965 10
D34965 N34965 0 diode
R34966 N34965 N34966 10
D34966 N34966 0 diode
R34967 N34966 N34967 10
D34967 N34967 0 diode
R34968 N34967 N34968 10
D34968 N34968 0 diode
R34969 N34968 N34969 10
D34969 N34969 0 diode
R34970 N34969 N34970 10
D34970 N34970 0 diode
R34971 N34970 N34971 10
D34971 N34971 0 diode
R34972 N34971 N34972 10
D34972 N34972 0 diode
R34973 N34972 N34973 10
D34973 N34973 0 diode
R34974 N34973 N34974 10
D34974 N34974 0 diode
R34975 N34974 N34975 10
D34975 N34975 0 diode
R34976 N34975 N34976 10
D34976 N34976 0 diode
R34977 N34976 N34977 10
D34977 N34977 0 diode
R34978 N34977 N34978 10
D34978 N34978 0 diode
R34979 N34978 N34979 10
D34979 N34979 0 diode
R34980 N34979 N34980 10
D34980 N34980 0 diode
R34981 N34980 N34981 10
D34981 N34981 0 diode
R34982 N34981 N34982 10
D34982 N34982 0 diode
R34983 N34982 N34983 10
D34983 N34983 0 diode
R34984 N34983 N34984 10
D34984 N34984 0 diode
R34985 N34984 N34985 10
D34985 N34985 0 diode
R34986 N34985 N34986 10
D34986 N34986 0 diode
R34987 N34986 N34987 10
D34987 N34987 0 diode
R34988 N34987 N34988 10
D34988 N34988 0 diode
R34989 N34988 N34989 10
D34989 N34989 0 diode
R34990 N34989 N34990 10
D34990 N34990 0 diode
R34991 N34990 N34991 10
D34991 N34991 0 diode
R34992 N34991 N34992 10
D34992 N34992 0 diode
R34993 N34992 N34993 10
D34993 N34993 0 diode
R34994 N34993 N34994 10
D34994 N34994 0 diode
R34995 N34994 N34995 10
D34995 N34995 0 diode
R34996 N34995 N34996 10
D34996 N34996 0 diode
R34997 N34996 N34997 10
D34997 N34997 0 diode
R34998 N34997 N34998 10
D34998 N34998 0 diode
R34999 N34998 N34999 10
D34999 N34999 0 diode
R35000 N34999 N35000 10
D35000 N35000 0 diode
R35001 N35000 N35001 10
D35001 N35001 0 diode
R35002 N35001 N35002 10
D35002 N35002 0 diode
R35003 N35002 N35003 10
D35003 N35003 0 diode
R35004 N35003 N35004 10
D35004 N35004 0 diode
R35005 N35004 N35005 10
D35005 N35005 0 diode
R35006 N35005 N35006 10
D35006 N35006 0 diode
R35007 N35006 N35007 10
D35007 N35007 0 diode
R35008 N35007 N35008 10
D35008 N35008 0 diode
R35009 N35008 N35009 10
D35009 N35009 0 diode
R35010 N35009 N35010 10
D35010 N35010 0 diode
R35011 N35010 N35011 10
D35011 N35011 0 diode
R35012 N35011 N35012 10
D35012 N35012 0 diode
R35013 N35012 N35013 10
D35013 N35013 0 diode
R35014 N35013 N35014 10
D35014 N35014 0 diode
R35015 N35014 N35015 10
D35015 N35015 0 diode
R35016 N35015 N35016 10
D35016 N35016 0 diode
R35017 N35016 N35017 10
D35017 N35017 0 diode
R35018 N35017 N35018 10
D35018 N35018 0 diode
R35019 N35018 N35019 10
D35019 N35019 0 diode
R35020 N35019 N35020 10
D35020 N35020 0 diode
R35021 N35020 N35021 10
D35021 N35021 0 diode
R35022 N35021 N35022 10
D35022 N35022 0 diode
R35023 N35022 N35023 10
D35023 N35023 0 diode
R35024 N35023 N35024 10
D35024 N35024 0 diode
R35025 N35024 N35025 10
D35025 N35025 0 diode
R35026 N35025 N35026 10
D35026 N35026 0 diode
R35027 N35026 N35027 10
D35027 N35027 0 diode
R35028 N35027 N35028 10
D35028 N35028 0 diode
R35029 N35028 N35029 10
D35029 N35029 0 diode
R35030 N35029 N35030 10
D35030 N35030 0 diode
R35031 N35030 N35031 10
D35031 N35031 0 diode
R35032 N35031 N35032 10
D35032 N35032 0 diode
R35033 N35032 N35033 10
D35033 N35033 0 diode
R35034 N35033 N35034 10
D35034 N35034 0 diode
R35035 N35034 N35035 10
D35035 N35035 0 diode
R35036 N35035 N35036 10
D35036 N35036 0 diode
R35037 N35036 N35037 10
D35037 N35037 0 diode
R35038 N35037 N35038 10
D35038 N35038 0 diode
R35039 N35038 N35039 10
D35039 N35039 0 diode
R35040 N35039 N35040 10
D35040 N35040 0 diode
R35041 N35040 N35041 10
D35041 N35041 0 diode
R35042 N35041 N35042 10
D35042 N35042 0 diode
R35043 N35042 N35043 10
D35043 N35043 0 diode
R35044 N35043 N35044 10
D35044 N35044 0 diode
R35045 N35044 N35045 10
D35045 N35045 0 diode
R35046 N35045 N35046 10
D35046 N35046 0 diode
R35047 N35046 N35047 10
D35047 N35047 0 diode
R35048 N35047 N35048 10
D35048 N35048 0 diode
R35049 N35048 N35049 10
D35049 N35049 0 diode
R35050 N35049 N35050 10
D35050 N35050 0 diode
R35051 N35050 N35051 10
D35051 N35051 0 diode
R35052 N35051 N35052 10
D35052 N35052 0 diode
R35053 N35052 N35053 10
D35053 N35053 0 diode
R35054 N35053 N35054 10
D35054 N35054 0 diode
R35055 N35054 N35055 10
D35055 N35055 0 diode
R35056 N35055 N35056 10
D35056 N35056 0 diode
R35057 N35056 N35057 10
D35057 N35057 0 diode
R35058 N35057 N35058 10
D35058 N35058 0 diode
R35059 N35058 N35059 10
D35059 N35059 0 diode
R35060 N35059 N35060 10
D35060 N35060 0 diode
R35061 N35060 N35061 10
D35061 N35061 0 diode
R35062 N35061 N35062 10
D35062 N35062 0 diode
R35063 N35062 N35063 10
D35063 N35063 0 diode
R35064 N35063 N35064 10
D35064 N35064 0 diode
R35065 N35064 N35065 10
D35065 N35065 0 diode
R35066 N35065 N35066 10
D35066 N35066 0 diode
R35067 N35066 N35067 10
D35067 N35067 0 diode
R35068 N35067 N35068 10
D35068 N35068 0 diode
R35069 N35068 N35069 10
D35069 N35069 0 diode
R35070 N35069 N35070 10
D35070 N35070 0 diode
R35071 N35070 N35071 10
D35071 N35071 0 diode
R35072 N35071 N35072 10
D35072 N35072 0 diode
R35073 N35072 N35073 10
D35073 N35073 0 diode
R35074 N35073 N35074 10
D35074 N35074 0 diode
R35075 N35074 N35075 10
D35075 N35075 0 diode
R35076 N35075 N35076 10
D35076 N35076 0 diode
R35077 N35076 N35077 10
D35077 N35077 0 diode
R35078 N35077 N35078 10
D35078 N35078 0 diode
R35079 N35078 N35079 10
D35079 N35079 0 diode
R35080 N35079 N35080 10
D35080 N35080 0 diode
R35081 N35080 N35081 10
D35081 N35081 0 diode
R35082 N35081 N35082 10
D35082 N35082 0 diode
R35083 N35082 N35083 10
D35083 N35083 0 diode
R35084 N35083 N35084 10
D35084 N35084 0 diode
R35085 N35084 N35085 10
D35085 N35085 0 diode
R35086 N35085 N35086 10
D35086 N35086 0 diode
R35087 N35086 N35087 10
D35087 N35087 0 diode
R35088 N35087 N35088 10
D35088 N35088 0 diode
R35089 N35088 N35089 10
D35089 N35089 0 diode
R35090 N35089 N35090 10
D35090 N35090 0 diode
R35091 N35090 N35091 10
D35091 N35091 0 diode
R35092 N35091 N35092 10
D35092 N35092 0 diode
R35093 N35092 N35093 10
D35093 N35093 0 diode
R35094 N35093 N35094 10
D35094 N35094 0 diode
R35095 N35094 N35095 10
D35095 N35095 0 diode
R35096 N35095 N35096 10
D35096 N35096 0 diode
R35097 N35096 N35097 10
D35097 N35097 0 diode
R35098 N35097 N35098 10
D35098 N35098 0 diode
R35099 N35098 N35099 10
D35099 N35099 0 diode
R35100 N35099 N35100 10
D35100 N35100 0 diode
R35101 N35100 N35101 10
D35101 N35101 0 diode
R35102 N35101 N35102 10
D35102 N35102 0 diode
R35103 N35102 N35103 10
D35103 N35103 0 diode
R35104 N35103 N35104 10
D35104 N35104 0 diode
R35105 N35104 N35105 10
D35105 N35105 0 diode
R35106 N35105 N35106 10
D35106 N35106 0 diode
R35107 N35106 N35107 10
D35107 N35107 0 diode
R35108 N35107 N35108 10
D35108 N35108 0 diode
R35109 N35108 N35109 10
D35109 N35109 0 diode
R35110 N35109 N35110 10
D35110 N35110 0 diode
R35111 N35110 N35111 10
D35111 N35111 0 diode
R35112 N35111 N35112 10
D35112 N35112 0 diode
R35113 N35112 N35113 10
D35113 N35113 0 diode
R35114 N35113 N35114 10
D35114 N35114 0 diode
R35115 N35114 N35115 10
D35115 N35115 0 diode
R35116 N35115 N35116 10
D35116 N35116 0 diode
R35117 N35116 N35117 10
D35117 N35117 0 diode
R35118 N35117 N35118 10
D35118 N35118 0 diode
R35119 N35118 N35119 10
D35119 N35119 0 diode
R35120 N35119 N35120 10
D35120 N35120 0 diode
R35121 N35120 N35121 10
D35121 N35121 0 diode
R35122 N35121 N35122 10
D35122 N35122 0 diode
R35123 N35122 N35123 10
D35123 N35123 0 diode
R35124 N35123 N35124 10
D35124 N35124 0 diode
R35125 N35124 N35125 10
D35125 N35125 0 diode
R35126 N35125 N35126 10
D35126 N35126 0 diode
R35127 N35126 N35127 10
D35127 N35127 0 diode
R35128 N35127 N35128 10
D35128 N35128 0 diode
R35129 N35128 N35129 10
D35129 N35129 0 diode
R35130 N35129 N35130 10
D35130 N35130 0 diode
R35131 N35130 N35131 10
D35131 N35131 0 diode
R35132 N35131 N35132 10
D35132 N35132 0 diode
R35133 N35132 N35133 10
D35133 N35133 0 diode
R35134 N35133 N35134 10
D35134 N35134 0 diode
R35135 N35134 N35135 10
D35135 N35135 0 diode
R35136 N35135 N35136 10
D35136 N35136 0 diode
R35137 N35136 N35137 10
D35137 N35137 0 diode
R35138 N35137 N35138 10
D35138 N35138 0 diode
R35139 N35138 N35139 10
D35139 N35139 0 diode
R35140 N35139 N35140 10
D35140 N35140 0 diode
R35141 N35140 N35141 10
D35141 N35141 0 diode
R35142 N35141 N35142 10
D35142 N35142 0 diode
R35143 N35142 N35143 10
D35143 N35143 0 diode
R35144 N35143 N35144 10
D35144 N35144 0 diode
R35145 N35144 N35145 10
D35145 N35145 0 diode
R35146 N35145 N35146 10
D35146 N35146 0 diode
R35147 N35146 N35147 10
D35147 N35147 0 diode
R35148 N35147 N35148 10
D35148 N35148 0 diode
R35149 N35148 N35149 10
D35149 N35149 0 diode
R35150 N35149 N35150 10
D35150 N35150 0 diode
R35151 N35150 N35151 10
D35151 N35151 0 diode
R35152 N35151 N35152 10
D35152 N35152 0 diode
R35153 N35152 N35153 10
D35153 N35153 0 diode
R35154 N35153 N35154 10
D35154 N35154 0 diode
R35155 N35154 N35155 10
D35155 N35155 0 diode
R35156 N35155 N35156 10
D35156 N35156 0 diode
R35157 N35156 N35157 10
D35157 N35157 0 diode
R35158 N35157 N35158 10
D35158 N35158 0 diode
R35159 N35158 N35159 10
D35159 N35159 0 diode
R35160 N35159 N35160 10
D35160 N35160 0 diode
R35161 N35160 N35161 10
D35161 N35161 0 diode
R35162 N35161 N35162 10
D35162 N35162 0 diode
R35163 N35162 N35163 10
D35163 N35163 0 diode
R35164 N35163 N35164 10
D35164 N35164 0 diode
R35165 N35164 N35165 10
D35165 N35165 0 diode
R35166 N35165 N35166 10
D35166 N35166 0 diode
R35167 N35166 N35167 10
D35167 N35167 0 diode
R35168 N35167 N35168 10
D35168 N35168 0 diode
R35169 N35168 N35169 10
D35169 N35169 0 diode
R35170 N35169 N35170 10
D35170 N35170 0 diode
R35171 N35170 N35171 10
D35171 N35171 0 diode
R35172 N35171 N35172 10
D35172 N35172 0 diode
R35173 N35172 N35173 10
D35173 N35173 0 diode
R35174 N35173 N35174 10
D35174 N35174 0 diode
R35175 N35174 N35175 10
D35175 N35175 0 diode
R35176 N35175 N35176 10
D35176 N35176 0 diode
R35177 N35176 N35177 10
D35177 N35177 0 diode
R35178 N35177 N35178 10
D35178 N35178 0 diode
R35179 N35178 N35179 10
D35179 N35179 0 diode
R35180 N35179 N35180 10
D35180 N35180 0 diode
R35181 N35180 N35181 10
D35181 N35181 0 diode
R35182 N35181 N35182 10
D35182 N35182 0 diode
R35183 N35182 N35183 10
D35183 N35183 0 diode
R35184 N35183 N35184 10
D35184 N35184 0 diode
R35185 N35184 N35185 10
D35185 N35185 0 diode
R35186 N35185 N35186 10
D35186 N35186 0 diode
R35187 N35186 N35187 10
D35187 N35187 0 diode
R35188 N35187 N35188 10
D35188 N35188 0 diode
R35189 N35188 N35189 10
D35189 N35189 0 diode
R35190 N35189 N35190 10
D35190 N35190 0 diode
R35191 N35190 N35191 10
D35191 N35191 0 diode
R35192 N35191 N35192 10
D35192 N35192 0 diode
R35193 N35192 N35193 10
D35193 N35193 0 diode
R35194 N35193 N35194 10
D35194 N35194 0 diode
R35195 N35194 N35195 10
D35195 N35195 0 diode
R35196 N35195 N35196 10
D35196 N35196 0 diode
R35197 N35196 N35197 10
D35197 N35197 0 diode
R35198 N35197 N35198 10
D35198 N35198 0 diode
R35199 N35198 N35199 10
D35199 N35199 0 diode
R35200 N35199 N35200 10
D35200 N35200 0 diode
R35201 N35200 N35201 10
D35201 N35201 0 diode
R35202 N35201 N35202 10
D35202 N35202 0 diode
R35203 N35202 N35203 10
D35203 N35203 0 diode
R35204 N35203 N35204 10
D35204 N35204 0 diode
R35205 N35204 N35205 10
D35205 N35205 0 diode
R35206 N35205 N35206 10
D35206 N35206 0 diode
R35207 N35206 N35207 10
D35207 N35207 0 diode
R35208 N35207 N35208 10
D35208 N35208 0 diode
R35209 N35208 N35209 10
D35209 N35209 0 diode
R35210 N35209 N35210 10
D35210 N35210 0 diode
R35211 N35210 N35211 10
D35211 N35211 0 diode
R35212 N35211 N35212 10
D35212 N35212 0 diode
R35213 N35212 N35213 10
D35213 N35213 0 diode
R35214 N35213 N35214 10
D35214 N35214 0 diode
R35215 N35214 N35215 10
D35215 N35215 0 diode
R35216 N35215 N35216 10
D35216 N35216 0 diode
R35217 N35216 N35217 10
D35217 N35217 0 diode
R35218 N35217 N35218 10
D35218 N35218 0 diode
R35219 N35218 N35219 10
D35219 N35219 0 diode
R35220 N35219 N35220 10
D35220 N35220 0 diode
R35221 N35220 N35221 10
D35221 N35221 0 diode
R35222 N35221 N35222 10
D35222 N35222 0 diode
R35223 N35222 N35223 10
D35223 N35223 0 diode
R35224 N35223 N35224 10
D35224 N35224 0 diode
R35225 N35224 N35225 10
D35225 N35225 0 diode
R35226 N35225 N35226 10
D35226 N35226 0 diode
R35227 N35226 N35227 10
D35227 N35227 0 diode
R35228 N35227 N35228 10
D35228 N35228 0 diode
R35229 N35228 N35229 10
D35229 N35229 0 diode
R35230 N35229 N35230 10
D35230 N35230 0 diode
R35231 N35230 N35231 10
D35231 N35231 0 diode
R35232 N35231 N35232 10
D35232 N35232 0 diode
R35233 N35232 N35233 10
D35233 N35233 0 diode
R35234 N35233 N35234 10
D35234 N35234 0 diode
R35235 N35234 N35235 10
D35235 N35235 0 diode
R35236 N35235 N35236 10
D35236 N35236 0 diode
R35237 N35236 N35237 10
D35237 N35237 0 diode
R35238 N35237 N35238 10
D35238 N35238 0 diode
R35239 N35238 N35239 10
D35239 N35239 0 diode
R35240 N35239 N35240 10
D35240 N35240 0 diode
R35241 N35240 N35241 10
D35241 N35241 0 diode
R35242 N35241 N35242 10
D35242 N35242 0 diode
R35243 N35242 N35243 10
D35243 N35243 0 diode
R35244 N35243 N35244 10
D35244 N35244 0 diode
R35245 N35244 N35245 10
D35245 N35245 0 diode
R35246 N35245 N35246 10
D35246 N35246 0 diode
R35247 N35246 N35247 10
D35247 N35247 0 diode
R35248 N35247 N35248 10
D35248 N35248 0 diode
R35249 N35248 N35249 10
D35249 N35249 0 diode
R35250 N35249 N35250 10
D35250 N35250 0 diode
R35251 N35250 N35251 10
D35251 N35251 0 diode
R35252 N35251 N35252 10
D35252 N35252 0 diode
R35253 N35252 N35253 10
D35253 N35253 0 diode
R35254 N35253 N35254 10
D35254 N35254 0 diode
R35255 N35254 N35255 10
D35255 N35255 0 diode
R35256 N35255 N35256 10
D35256 N35256 0 diode
R35257 N35256 N35257 10
D35257 N35257 0 diode
R35258 N35257 N35258 10
D35258 N35258 0 diode
R35259 N35258 N35259 10
D35259 N35259 0 diode
R35260 N35259 N35260 10
D35260 N35260 0 diode
R35261 N35260 N35261 10
D35261 N35261 0 diode
R35262 N35261 N35262 10
D35262 N35262 0 diode
R35263 N35262 N35263 10
D35263 N35263 0 diode
R35264 N35263 N35264 10
D35264 N35264 0 diode
R35265 N35264 N35265 10
D35265 N35265 0 diode
R35266 N35265 N35266 10
D35266 N35266 0 diode
R35267 N35266 N35267 10
D35267 N35267 0 diode
R35268 N35267 N35268 10
D35268 N35268 0 diode
R35269 N35268 N35269 10
D35269 N35269 0 diode
R35270 N35269 N35270 10
D35270 N35270 0 diode
R35271 N35270 N35271 10
D35271 N35271 0 diode
R35272 N35271 N35272 10
D35272 N35272 0 diode
R35273 N35272 N35273 10
D35273 N35273 0 diode
R35274 N35273 N35274 10
D35274 N35274 0 diode
R35275 N35274 N35275 10
D35275 N35275 0 diode
R35276 N35275 N35276 10
D35276 N35276 0 diode
R35277 N35276 N35277 10
D35277 N35277 0 diode
R35278 N35277 N35278 10
D35278 N35278 0 diode
R35279 N35278 N35279 10
D35279 N35279 0 diode
R35280 N35279 N35280 10
D35280 N35280 0 diode
R35281 N35280 N35281 10
D35281 N35281 0 diode
R35282 N35281 N35282 10
D35282 N35282 0 diode
R35283 N35282 N35283 10
D35283 N35283 0 diode
R35284 N35283 N35284 10
D35284 N35284 0 diode
R35285 N35284 N35285 10
D35285 N35285 0 diode
R35286 N35285 N35286 10
D35286 N35286 0 diode
R35287 N35286 N35287 10
D35287 N35287 0 diode
R35288 N35287 N35288 10
D35288 N35288 0 diode
R35289 N35288 N35289 10
D35289 N35289 0 diode
R35290 N35289 N35290 10
D35290 N35290 0 diode
R35291 N35290 N35291 10
D35291 N35291 0 diode
R35292 N35291 N35292 10
D35292 N35292 0 diode
R35293 N35292 N35293 10
D35293 N35293 0 diode
R35294 N35293 N35294 10
D35294 N35294 0 diode
R35295 N35294 N35295 10
D35295 N35295 0 diode
R35296 N35295 N35296 10
D35296 N35296 0 diode
R35297 N35296 N35297 10
D35297 N35297 0 diode
R35298 N35297 N35298 10
D35298 N35298 0 diode
R35299 N35298 N35299 10
D35299 N35299 0 diode
R35300 N35299 N35300 10
D35300 N35300 0 diode
R35301 N35300 N35301 10
D35301 N35301 0 diode
R35302 N35301 N35302 10
D35302 N35302 0 diode
R35303 N35302 N35303 10
D35303 N35303 0 diode
R35304 N35303 N35304 10
D35304 N35304 0 diode
R35305 N35304 N35305 10
D35305 N35305 0 diode
R35306 N35305 N35306 10
D35306 N35306 0 diode
R35307 N35306 N35307 10
D35307 N35307 0 diode
R35308 N35307 N35308 10
D35308 N35308 0 diode
R35309 N35308 N35309 10
D35309 N35309 0 diode
R35310 N35309 N35310 10
D35310 N35310 0 diode
R35311 N35310 N35311 10
D35311 N35311 0 diode
R35312 N35311 N35312 10
D35312 N35312 0 diode
R35313 N35312 N35313 10
D35313 N35313 0 diode
R35314 N35313 N35314 10
D35314 N35314 0 diode
R35315 N35314 N35315 10
D35315 N35315 0 diode
R35316 N35315 N35316 10
D35316 N35316 0 diode
R35317 N35316 N35317 10
D35317 N35317 0 diode
R35318 N35317 N35318 10
D35318 N35318 0 diode
R35319 N35318 N35319 10
D35319 N35319 0 diode
R35320 N35319 N35320 10
D35320 N35320 0 diode
R35321 N35320 N35321 10
D35321 N35321 0 diode
R35322 N35321 N35322 10
D35322 N35322 0 diode
R35323 N35322 N35323 10
D35323 N35323 0 diode
R35324 N35323 N35324 10
D35324 N35324 0 diode
R35325 N35324 N35325 10
D35325 N35325 0 diode
R35326 N35325 N35326 10
D35326 N35326 0 diode
R35327 N35326 N35327 10
D35327 N35327 0 diode
R35328 N35327 N35328 10
D35328 N35328 0 diode
R35329 N35328 N35329 10
D35329 N35329 0 diode
R35330 N35329 N35330 10
D35330 N35330 0 diode
R35331 N35330 N35331 10
D35331 N35331 0 diode
R35332 N35331 N35332 10
D35332 N35332 0 diode
R35333 N35332 N35333 10
D35333 N35333 0 diode
R35334 N35333 N35334 10
D35334 N35334 0 diode
R35335 N35334 N35335 10
D35335 N35335 0 diode
R35336 N35335 N35336 10
D35336 N35336 0 diode
R35337 N35336 N35337 10
D35337 N35337 0 diode
R35338 N35337 N35338 10
D35338 N35338 0 diode
R35339 N35338 N35339 10
D35339 N35339 0 diode
R35340 N35339 N35340 10
D35340 N35340 0 diode
R35341 N35340 N35341 10
D35341 N35341 0 diode
R35342 N35341 N35342 10
D35342 N35342 0 diode
R35343 N35342 N35343 10
D35343 N35343 0 diode
R35344 N35343 N35344 10
D35344 N35344 0 diode
R35345 N35344 N35345 10
D35345 N35345 0 diode
R35346 N35345 N35346 10
D35346 N35346 0 diode
R35347 N35346 N35347 10
D35347 N35347 0 diode
R35348 N35347 N35348 10
D35348 N35348 0 diode
R35349 N35348 N35349 10
D35349 N35349 0 diode
R35350 N35349 N35350 10
D35350 N35350 0 diode
R35351 N35350 N35351 10
D35351 N35351 0 diode
R35352 N35351 N35352 10
D35352 N35352 0 diode
R35353 N35352 N35353 10
D35353 N35353 0 diode
R35354 N35353 N35354 10
D35354 N35354 0 diode
R35355 N35354 N35355 10
D35355 N35355 0 diode
R35356 N35355 N35356 10
D35356 N35356 0 diode
R35357 N35356 N35357 10
D35357 N35357 0 diode
R35358 N35357 N35358 10
D35358 N35358 0 diode
R35359 N35358 N35359 10
D35359 N35359 0 diode
R35360 N35359 N35360 10
D35360 N35360 0 diode
R35361 N35360 N35361 10
D35361 N35361 0 diode
R35362 N35361 N35362 10
D35362 N35362 0 diode
R35363 N35362 N35363 10
D35363 N35363 0 diode
R35364 N35363 N35364 10
D35364 N35364 0 diode
R35365 N35364 N35365 10
D35365 N35365 0 diode
R35366 N35365 N35366 10
D35366 N35366 0 diode
R35367 N35366 N35367 10
D35367 N35367 0 diode
R35368 N35367 N35368 10
D35368 N35368 0 diode
R35369 N35368 N35369 10
D35369 N35369 0 diode
R35370 N35369 N35370 10
D35370 N35370 0 diode
R35371 N35370 N35371 10
D35371 N35371 0 diode
R35372 N35371 N35372 10
D35372 N35372 0 diode
R35373 N35372 N35373 10
D35373 N35373 0 diode
R35374 N35373 N35374 10
D35374 N35374 0 diode
R35375 N35374 N35375 10
D35375 N35375 0 diode
R35376 N35375 N35376 10
D35376 N35376 0 diode
R35377 N35376 N35377 10
D35377 N35377 0 diode
R35378 N35377 N35378 10
D35378 N35378 0 diode
R35379 N35378 N35379 10
D35379 N35379 0 diode
R35380 N35379 N35380 10
D35380 N35380 0 diode
R35381 N35380 N35381 10
D35381 N35381 0 diode
R35382 N35381 N35382 10
D35382 N35382 0 diode
R35383 N35382 N35383 10
D35383 N35383 0 diode
R35384 N35383 N35384 10
D35384 N35384 0 diode
R35385 N35384 N35385 10
D35385 N35385 0 diode
R35386 N35385 N35386 10
D35386 N35386 0 diode
R35387 N35386 N35387 10
D35387 N35387 0 diode
R35388 N35387 N35388 10
D35388 N35388 0 diode
R35389 N35388 N35389 10
D35389 N35389 0 diode
R35390 N35389 N35390 10
D35390 N35390 0 diode
R35391 N35390 N35391 10
D35391 N35391 0 diode
R35392 N35391 N35392 10
D35392 N35392 0 diode
R35393 N35392 N35393 10
D35393 N35393 0 diode
R35394 N35393 N35394 10
D35394 N35394 0 diode
R35395 N35394 N35395 10
D35395 N35395 0 diode
R35396 N35395 N35396 10
D35396 N35396 0 diode
R35397 N35396 N35397 10
D35397 N35397 0 diode
R35398 N35397 N35398 10
D35398 N35398 0 diode
R35399 N35398 N35399 10
D35399 N35399 0 diode
R35400 N35399 N35400 10
D35400 N35400 0 diode
R35401 N35400 N35401 10
D35401 N35401 0 diode
R35402 N35401 N35402 10
D35402 N35402 0 diode
R35403 N35402 N35403 10
D35403 N35403 0 diode
R35404 N35403 N35404 10
D35404 N35404 0 diode
R35405 N35404 N35405 10
D35405 N35405 0 diode
R35406 N35405 N35406 10
D35406 N35406 0 diode
R35407 N35406 N35407 10
D35407 N35407 0 diode
R35408 N35407 N35408 10
D35408 N35408 0 diode
R35409 N35408 N35409 10
D35409 N35409 0 diode
R35410 N35409 N35410 10
D35410 N35410 0 diode
R35411 N35410 N35411 10
D35411 N35411 0 diode
R35412 N35411 N35412 10
D35412 N35412 0 diode
R35413 N35412 N35413 10
D35413 N35413 0 diode
R35414 N35413 N35414 10
D35414 N35414 0 diode
R35415 N35414 N35415 10
D35415 N35415 0 diode
R35416 N35415 N35416 10
D35416 N35416 0 diode
R35417 N35416 N35417 10
D35417 N35417 0 diode
R35418 N35417 N35418 10
D35418 N35418 0 diode
R35419 N35418 N35419 10
D35419 N35419 0 diode
R35420 N35419 N35420 10
D35420 N35420 0 diode
R35421 N35420 N35421 10
D35421 N35421 0 diode
R35422 N35421 N35422 10
D35422 N35422 0 diode
R35423 N35422 N35423 10
D35423 N35423 0 diode
R35424 N35423 N35424 10
D35424 N35424 0 diode
R35425 N35424 N35425 10
D35425 N35425 0 diode
R35426 N35425 N35426 10
D35426 N35426 0 diode
R35427 N35426 N35427 10
D35427 N35427 0 diode
R35428 N35427 N35428 10
D35428 N35428 0 diode
R35429 N35428 N35429 10
D35429 N35429 0 diode
R35430 N35429 N35430 10
D35430 N35430 0 diode
R35431 N35430 N35431 10
D35431 N35431 0 diode
R35432 N35431 N35432 10
D35432 N35432 0 diode
R35433 N35432 N35433 10
D35433 N35433 0 diode
R35434 N35433 N35434 10
D35434 N35434 0 diode
R35435 N35434 N35435 10
D35435 N35435 0 diode
R35436 N35435 N35436 10
D35436 N35436 0 diode
R35437 N35436 N35437 10
D35437 N35437 0 diode
R35438 N35437 N35438 10
D35438 N35438 0 diode
R35439 N35438 N35439 10
D35439 N35439 0 diode
R35440 N35439 N35440 10
D35440 N35440 0 diode
R35441 N35440 N35441 10
D35441 N35441 0 diode
R35442 N35441 N35442 10
D35442 N35442 0 diode
R35443 N35442 N35443 10
D35443 N35443 0 diode
R35444 N35443 N35444 10
D35444 N35444 0 diode
R35445 N35444 N35445 10
D35445 N35445 0 diode
R35446 N35445 N35446 10
D35446 N35446 0 diode
R35447 N35446 N35447 10
D35447 N35447 0 diode
R35448 N35447 N35448 10
D35448 N35448 0 diode
R35449 N35448 N35449 10
D35449 N35449 0 diode
R35450 N35449 N35450 10
D35450 N35450 0 diode
R35451 N35450 N35451 10
D35451 N35451 0 diode
R35452 N35451 N35452 10
D35452 N35452 0 diode
R35453 N35452 N35453 10
D35453 N35453 0 diode
R35454 N35453 N35454 10
D35454 N35454 0 diode
R35455 N35454 N35455 10
D35455 N35455 0 diode
R35456 N35455 N35456 10
D35456 N35456 0 diode
R35457 N35456 N35457 10
D35457 N35457 0 diode
R35458 N35457 N35458 10
D35458 N35458 0 diode
R35459 N35458 N35459 10
D35459 N35459 0 diode
R35460 N35459 N35460 10
D35460 N35460 0 diode
R35461 N35460 N35461 10
D35461 N35461 0 diode
R35462 N35461 N35462 10
D35462 N35462 0 diode
R35463 N35462 N35463 10
D35463 N35463 0 diode
R35464 N35463 N35464 10
D35464 N35464 0 diode
R35465 N35464 N35465 10
D35465 N35465 0 diode
R35466 N35465 N35466 10
D35466 N35466 0 diode
R35467 N35466 N35467 10
D35467 N35467 0 diode
R35468 N35467 N35468 10
D35468 N35468 0 diode
R35469 N35468 N35469 10
D35469 N35469 0 diode
R35470 N35469 N35470 10
D35470 N35470 0 diode
R35471 N35470 N35471 10
D35471 N35471 0 diode
R35472 N35471 N35472 10
D35472 N35472 0 diode
R35473 N35472 N35473 10
D35473 N35473 0 diode
R35474 N35473 N35474 10
D35474 N35474 0 diode
R35475 N35474 N35475 10
D35475 N35475 0 diode
R35476 N35475 N35476 10
D35476 N35476 0 diode
R35477 N35476 N35477 10
D35477 N35477 0 diode
R35478 N35477 N35478 10
D35478 N35478 0 diode
R35479 N35478 N35479 10
D35479 N35479 0 diode
R35480 N35479 N35480 10
D35480 N35480 0 diode
R35481 N35480 N35481 10
D35481 N35481 0 diode
R35482 N35481 N35482 10
D35482 N35482 0 diode
R35483 N35482 N35483 10
D35483 N35483 0 diode
R35484 N35483 N35484 10
D35484 N35484 0 diode
R35485 N35484 N35485 10
D35485 N35485 0 diode
R35486 N35485 N35486 10
D35486 N35486 0 diode
R35487 N35486 N35487 10
D35487 N35487 0 diode
R35488 N35487 N35488 10
D35488 N35488 0 diode
R35489 N35488 N35489 10
D35489 N35489 0 diode
R35490 N35489 N35490 10
D35490 N35490 0 diode
R35491 N35490 N35491 10
D35491 N35491 0 diode
R35492 N35491 N35492 10
D35492 N35492 0 diode
R35493 N35492 N35493 10
D35493 N35493 0 diode
R35494 N35493 N35494 10
D35494 N35494 0 diode
R35495 N35494 N35495 10
D35495 N35495 0 diode
R35496 N35495 N35496 10
D35496 N35496 0 diode
R35497 N35496 N35497 10
D35497 N35497 0 diode
R35498 N35497 N35498 10
D35498 N35498 0 diode
R35499 N35498 N35499 10
D35499 N35499 0 diode
R35500 N35499 N35500 10
D35500 N35500 0 diode
R35501 N35500 N35501 10
D35501 N35501 0 diode
R35502 N35501 N35502 10
D35502 N35502 0 diode
R35503 N35502 N35503 10
D35503 N35503 0 diode
R35504 N35503 N35504 10
D35504 N35504 0 diode
R35505 N35504 N35505 10
D35505 N35505 0 diode
R35506 N35505 N35506 10
D35506 N35506 0 diode
R35507 N35506 N35507 10
D35507 N35507 0 diode
R35508 N35507 N35508 10
D35508 N35508 0 diode
R35509 N35508 N35509 10
D35509 N35509 0 diode
R35510 N35509 N35510 10
D35510 N35510 0 diode
R35511 N35510 N35511 10
D35511 N35511 0 diode
R35512 N35511 N35512 10
D35512 N35512 0 diode
R35513 N35512 N35513 10
D35513 N35513 0 diode
R35514 N35513 N35514 10
D35514 N35514 0 diode
R35515 N35514 N35515 10
D35515 N35515 0 diode
R35516 N35515 N35516 10
D35516 N35516 0 diode
R35517 N35516 N35517 10
D35517 N35517 0 diode
R35518 N35517 N35518 10
D35518 N35518 0 diode
R35519 N35518 N35519 10
D35519 N35519 0 diode
R35520 N35519 N35520 10
D35520 N35520 0 diode
R35521 N35520 N35521 10
D35521 N35521 0 diode
R35522 N35521 N35522 10
D35522 N35522 0 diode
R35523 N35522 N35523 10
D35523 N35523 0 diode
R35524 N35523 N35524 10
D35524 N35524 0 diode
R35525 N35524 N35525 10
D35525 N35525 0 diode
R35526 N35525 N35526 10
D35526 N35526 0 diode
R35527 N35526 N35527 10
D35527 N35527 0 diode
R35528 N35527 N35528 10
D35528 N35528 0 diode
R35529 N35528 N35529 10
D35529 N35529 0 diode
R35530 N35529 N35530 10
D35530 N35530 0 diode
R35531 N35530 N35531 10
D35531 N35531 0 diode
R35532 N35531 N35532 10
D35532 N35532 0 diode
R35533 N35532 N35533 10
D35533 N35533 0 diode
R35534 N35533 N35534 10
D35534 N35534 0 diode
R35535 N35534 N35535 10
D35535 N35535 0 diode
R35536 N35535 N35536 10
D35536 N35536 0 diode
R35537 N35536 N35537 10
D35537 N35537 0 diode
R35538 N35537 N35538 10
D35538 N35538 0 diode
R35539 N35538 N35539 10
D35539 N35539 0 diode
R35540 N35539 N35540 10
D35540 N35540 0 diode
R35541 N35540 N35541 10
D35541 N35541 0 diode
R35542 N35541 N35542 10
D35542 N35542 0 diode
R35543 N35542 N35543 10
D35543 N35543 0 diode
R35544 N35543 N35544 10
D35544 N35544 0 diode
R35545 N35544 N35545 10
D35545 N35545 0 diode
R35546 N35545 N35546 10
D35546 N35546 0 diode
R35547 N35546 N35547 10
D35547 N35547 0 diode
R35548 N35547 N35548 10
D35548 N35548 0 diode
R35549 N35548 N35549 10
D35549 N35549 0 diode
R35550 N35549 N35550 10
D35550 N35550 0 diode
R35551 N35550 N35551 10
D35551 N35551 0 diode
R35552 N35551 N35552 10
D35552 N35552 0 diode
R35553 N35552 N35553 10
D35553 N35553 0 diode
R35554 N35553 N35554 10
D35554 N35554 0 diode
R35555 N35554 N35555 10
D35555 N35555 0 diode
R35556 N35555 N35556 10
D35556 N35556 0 diode
R35557 N35556 N35557 10
D35557 N35557 0 diode
R35558 N35557 N35558 10
D35558 N35558 0 diode
R35559 N35558 N35559 10
D35559 N35559 0 diode
R35560 N35559 N35560 10
D35560 N35560 0 diode
R35561 N35560 N35561 10
D35561 N35561 0 diode
R35562 N35561 N35562 10
D35562 N35562 0 diode
R35563 N35562 N35563 10
D35563 N35563 0 diode
R35564 N35563 N35564 10
D35564 N35564 0 diode
R35565 N35564 N35565 10
D35565 N35565 0 diode
R35566 N35565 N35566 10
D35566 N35566 0 diode
R35567 N35566 N35567 10
D35567 N35567 0 diode
R35568 N35567 N35568 10
D35568 N35568 0 diode
R35569 N35568 N35569 10
D35569 N35569 0 diode
R35570 N35569 N35570 10
D35570 N35570 0 diode
R35571 N35570 N35571 10
D35571 N35571 0 diode
R35572 N35571 N35572 10
D35572 N35572 0 diode
R35573 N35572 N35573 10
D35573 N35573 0 diode
R35574 N35573 N35574 10
D35574 N35574 0 diode
R35575 N35574 N35575 10
D35575 N35575 0 diode
R35576 N35575 N35576 10
D35576 N35576 0 diode
R35577 N35576 N35577 10
D35577 N35577 0 diode
R35578 N35577 N35578 10
D35578 N35578 0 diode
R35579 N35578 N35579 10
D35579 N35579 0 diode
R35580 N35579 N35580 10
D35580 N35580 0 diode
R35581 N35580 N35581 10
D35581 N35581 0 diode
R35582 N35581 N35582 10
D35582 N35582 0 diode
R35583 N35582 N35583 10
D35583 N35583 0 diode
R35584 N35583 N35584 10
D35584 N35584 0 diode
R35585 N35584 N35585 10
D35585 N35585 0 diode
R35586 N35585 N35586 10
D35586 N35586 0 diode
R35587 N35586 N35587 10
D35587 N35587 0 diode
R35588 N35587 N35588 10
D35588 N35588 0 diode
R35589 N35588 N35589 10
D35589 N35589 0 diode
R35590 N35589 N35590 10
D35590 N35590 0 diode
R35591 N35590 N35591 10
D35591 N35591 0 diode
R35592 N35591 N35592 10
D35592 N35592 0 diode
R35593 N35592 N35593 10
D35593 N35593 0 diode
R35594 N35593 N35594 10
D35594 N35594 0 diode
R35595 N35594 N35595 10
D35595 N35595 0 diode
R35596 N35595 N35596 10
D35596 N35596 0 diode
R35597 N35596 N35597 10
D35597 N35597 0 diode
R35598 N35597 N35598 10
D35598 N35598 0 diode
R35599 N35598 N35599 10
D35599 N35599 0 diode
R35600 N35599 N35600 10
D35600 N35600 0 diode
R35601 N35600 N35601 10
D35601 N35601 0 diode
R35602 N35601 N35602 10
D35602 N35602 0 diode
R35603 N35602 N35603 10
D35603 N35603 0 diode
R35604 N35603 N35604 10
D35604 N35604 0 diode
R35605 N35604 N35605 10
D35605 N35605 0 diode
R35606 N35605 N35606 10
D35606 N35606 0 diode
R35607 N35606 N35607 10
D35607 N35607 0 diode
R35608 N35607 N35608 10
D35608 N35608 0 diode
R35609 N35608 N35609 10
D35609 N35609 0 diode
R35610 N35609 N35610 10
D35610 N35610 0 diode
R35611 N35610 N35611 10
D35611 N35611 0 diode
R35612 N35611 N35612 10
D35612 N35612 0 diode
R35613 N35612 N35613 10
D35613 N35613 0 diode
R35614 N35613 N35614 10
D35614 N35614 0 diode
R35615 N35614 N35615 10
D35615 N35615 0 diode
R35616 N35615 N35616 10
D35616 N35616 0 diode
R35617 N35616 N35617 10
D35617 N35617 0 diode
R35618 N35617 N35618 10
D35618 N35618 0 diode
R35619 N35618 N35619 10
D35619 N35619 0 diode
R35620 N35619 N35620 10
D35620 N35620 0 diode
R35621 N35620 N35621 10
D35621 N35621 0 diode
R35622 N35621 N35622 10
D35622 N35622 0 diode
R35623 N35622 N35623 10
D35623 N35623 0 diode
R35624 N35623 N35624 10
D35624 N35624 0 diode
R35625 N35624 N35625 10
D35625 N35625 0 diode
R35626 N35625 N35626 10
D35626 N35626 0 diode
R35627 N35626 N35627 10
D35627 N35627 0 diode
R35628 N35627 N35628 10
D35628 N35628 0 diode
R35629 N35628 N35629 10
D35629 N35629 0 diode
R35630 N35629 N35630 10
D35630 N35630 0 diode
R35631 N35630 N35631 10
D35631 N35631 0 diode
R35632 N35631 N35632 10
D35632 N35632 0 diode
R35633 N35632 N35633 10
D35633 N35633 0 diode
R35634 N35633 N35634 10
D35634 N35634 0 diode
R35635 N35634 N35635 10
D35635 N35635 0 diode
R35636 N35635 N35636 10
D35636 N35636 0 diode
R35637 N35636 N35637 10
D35637 N35637 0 diode
R35638 N35637 N35638 10
D35638 N35638 0 diode
R35639 N35638 N35639 10
D35639 N35639 0 diode
R35640 N35639 N35640 10
D35640 N35640 0 diode
R35641 N35640 N35641 10
D35641 N35641 0 diode
R35642 N35641 N35642 10
D35642 N35642 0 diode
R35643 N35642 N35643 10
D35643 N35643 0 diode
R35644 N35643 N35644 10
D35644 N35644 0 diode
R35645 N35644 N35645 10
D35645 N35645 0 diode
R35646 N35645 N35646 10
D35646 N35646 0 diode
R35647 N35646 N35647 10
D35647 N35647 0 diode
R35648 N35647 N35648 10
D35648 N35648 0 diode
R35649 N35648 N35649 10
D35649 N35649 0 diode
R35650 N35649 N35650 10
D35650 N35650 0 diode
R35651 N35650 N35651 10
D35651 N35651 0 diode
R35652 N35651 N35652 10
D35652 N35652 0 diode
R35653 N35652 N35653 10
D35653 N35653 0 diode
R35654 N35653 N35654 10
D35654 N35654 0 diode
R35655 N35654 N35655 10
D35655 N35655 0 diode
R35656 N35655 N35656 10
D35656 N35656 0 diode
R35657 N35656 N35657 10
D35657 N35657 0 diode
R35658 N35657 N35658 10
D35658 N35658 0 diode
R35659 N35658 N35659 10
D35659 N35659 0 diode
R35660 N35659 N35660 10
D35660 N35660 0 diode
R35661 N35660 N35661 10
D35661 N35661 0 diode
R35662 N35661 N35662 10
D35662 N35662 0 diode
R35663 N35662 N35663 10
D35663 N35663 0 diode
R35664 N35663 N35664 10
D35664 N35664 0 diode
R35665 N35664 N35665 10
D35665 N35665 0 diode
R35666 N35665 N35666 10
D35666 N35666 0 diode
R35667 N35666 N35667 10
D35667 N35667 0 diode
R35668 N35667 N35668 10
D35668 N35668 0 diode
R35669 N35668 N35669 10
D35669 N35669 0 diode
R35670 N35669 N35670 10
D35670 N35670 0 diode
R35671 N35670 N35671 10
D35671 N35671 0 diode
R35672 N35671 N35672 10
D35672 N35672 0 diode
R35673 N35672 N35673 10
D35673 N35673 0 diode
R35674 N35673 N35674 10
D35674 N35674 0 diode
R35675 N35674 N35675 10
D35675 N35675 0 diode
R35676 N35675 N35676 10
D35676 N35676 0 diode
R35677 N35676 N35677 10
D35677 N35677 0 diode
R35678 N35677 N35678 10
D35678 N35678 0 diode
R35679 N35678 N35679 10
D35679 N35679 0 diode
R35680 N35679 N35680 10
D35680 N35680 0 diode
R35681 N35680 N35681 10
D35681 N35681 0 diode
R35682 N35681 N35682 10
D35682 N35682 0 diode
R35683 N35682 N35683 10
D35683 N35683 0 diode
R35684 N35683 N35684 10
D35684 N35684 0 diode
R35685 N35684 N35685 10
D35685 N35685 0 diode
R35686 N35685 N35686 10
D35686 N35686 0 diode
R35687 N35686 N35687 10
D35687 N35687 0 diode
R35688 N35687 N35688 10
D35688 N35688 0 diode
R35689 N35688 N35689 10
D35689 N35689 0 diode
R35690 N35689 N35690 10
D35690 N35690 0 diode
R35691 N35690 N35691 10
D35691 N35691 0 diode
R35692 N35691 N35692 10
D35692 N35692 0 diode
R35693 N35692 N35693 10
D35693 N35693 0 diode
R35694 N35693 N35694 10
D35694 N35694 0 diode
R35695 N35694 N35695 10
D35695 N35695 0 diode
R35696 N35695 N35696 10
D35696 N35696 0 diode
R35697 N35696 N35697 10
D35697 N35697 0 diode
R35698 N35697 N35698 10
D35698 N35698 0 diode
R35699 N35698 N35699 10
D35699 N35699 0 diode
R35700 N35699 N35700 10
D35700 N35700 0 diode
R35701 N35700 N35701 10
D35701 N35701 0 diode
R35702 N35701 N35702 10
D35702 N35702 0 diode
R35703 N35702 N35703 10
D35703 N35703 0 diode
R35704 N35703 N35704 10
D35704 N35704 0 diode
R35705 N35704 N35705 10
D35705 N35705 0 diode
R35706 N35705 N35706 10
D35706 N35706 0 diode
R35707 N35706 N35707 10
D35707 N35707 0 diode
R35708 N35707 N35708 10
D35708 N35708 0 diode
R35709 N35708 N35709 10
D35709 N35709 0 diode
R35710 N35709 N35710 10
D35710 N35710 0 diode
R35711 N35710 N35711 10
D35711 N35711 0 diode
R35712 N35711 N35712 10
D35712 N35712 0 diode
R35713 N35712 N35713 10
D35713 N35713 0 diode
R35714 N35713 N35714 10
D35714 N35714 0 diode
R35715 N35714 N35715 10
D35715 N35715 0 diode
R35716 N35715 N35716 10
D35716 N35716 0 diode
R35717 N35716 N35717 10
D35717 N35717 0 diode
R35718 N35717 N35718 10
D35718 N35718 0 diode
R35719 N35718 N35719 10
D35719 N35719 0 diode
R35720 N35719 N35720 10
D35720 N35720 0 diode
R35721 N35720 N35721 10
D35721 N35721 0 diode
R35722 N35721 N35722 10
D35722 N35722 0 diode
R35723 N35722 N35723 10
D35723 N35723 0 diode
R35724 N35723 N35724 10
D35724 N35724 0 diode
R35725 N35724 N35725 10
D35725 N35725 0 diode
R35726 N35725 N35726 10
D35726 N35726 0 diode
R35727 N35726 N35727 10
D35727 N35727 0 diode
R35728 N35727 N35728 10
D35728 N35728 0 diode
R35729 N35728 N35729 10
D35729 N35729 0 diode
R35730 N35729 N35730 10
D35730 N35730 0 diode
R35731 N35730 N35731 10
D35731 N35731 0 diode
R35732 N35731 N35732 10
D35732 N35732 0 diode
R35733 N35732 N35733 10
D35733 N35733 0 diode
R35734 N35733 N35734 10
D35734 N35734 0 diode
R35735 N35734 N35735 10
D35735 N35735 0 diode
R35736 N35735 N35736 10
D35736 N35736 0 diode
R35737 N35736 N35737 10
D35737 N35737 0 diode
R35738 N35737 N35738 10
D35738 N35738 0 diode
R35739 N35738 N35739 10
D35739 N35739 0 diode
R35740 N35739 N35740 10
D35740 N35740 0 diode
R35741 N35740 N35741 10
D35741 N35741 0 diode
R35742 N35741 N35742 10
D35742 N35742 0 diode
R35743 N35742 N35743 10
D35743 N35743 0 diode
R35744 N35743 N35744 10
D35744 N35744 0 diode
R35745 N35744 N35745 10
D35745 N35745 0 diode
R35746 N35745 N35746 10
D35746 N35746 0 diode
R35747 N35746 N35747 10
D35747 N35747 0 diode
R35748 N35747 N35748 10
D35748 N35748 0 diode
R35749 N35748 N35749 10
D35749 N35749 0 diode
R35750 N35749 N35750 10
D35750 N35750 0 diode
R35751 N35750 N35751 10
D35751 N35751 0 diode
R35752 N35751 N35752 10
D35752 N35752 0 diode
R35753 N35752 N35753 10
D35753 N35753 0 diode
R35754 N35753 N35754 10
D35754 N35754 0 diode
R35755 N35754 N35755 10
D35755 N35755 0 diode
R35756 N35755 N35756 10
D35756 N35756 0 diode
R35757 N35756 N35757 10
D35757 N35757 0 diode
R35758 N35757 N35758 10
D35758 N35758 0 diode
R35759 N35758 N35759 10
D35759 N35759 0 diode
R35760 N35759 N35760 10
D35760 N35760 0 diode
R35761 N35760 N35761 10
D35761 N35761 0 diode
R35762 N35761 N35762 10
D35762 N35762 0 diode
R35763 N35762 N35763 10
D35763 N35763 0 diode
R35764 N35763 N35764 10
D35764 N35764 0 diode
R35765 N35764 N35765 10
D35765 N35765 0 diode
R35766 N35765 N35766 10
D35766 N35766 0 diode
R35767 N35766 N35767 10
D35767 N35767 0 diode
R35768 N35767 N35768 10
D35768 N35768 0 diode
R35769 N35768 N35769 10
D35769 N35769 0 diode
R35770 N35769 N35770 10
D35770 N35770 0 diode
R35771 N35770 N35771 10
D35771 N35771 0 diode
R35772 N35771 N35772 10
D35772 N35772 0 diode
R35773 N35772 N35773 10
D35773 N35773 0 diode
R35774 N35773 N35774 10
D35774 N35774 0 diode
R35775 N35774 N35775 10
D35775 N35775 0 diode
R35776 N35775 N35776 10
D35776 N35776 0 diode
R35777 N35776 N35777 10
D35777 N35777 0 diode
R35778 N35777 N35778 10
D35778 N35778 0 diode
R35779 N35778 N35779 10
D35779 N35779 0 diode
R35780 N35779 N35780 10
D35780 N35780 0 diode
R35781 N35780 N35781 10
D35781 N35781 0 diode
R35782 N35781 N35782 10
D35782 N35782 0 diode
R35783 N35782 N35783 10
D35783 N35783 0 diode
R35784 N35783 N35784 10
D35784 N35784 0 diode
R35785 N35784 N35785 10
D35785 N35785 0 diode
R35786 N35785 N35786 10
D35786 N35786 0 diode
R35787 N35786 N35787 10
D35787 N35787 0 diode
R35788 N35787 N35788 10
D35788 N35788 0 diode
R35789 N35788 N35789 10
D35789 N35789 0 diode
R35790 N35789 N35790 10
D35790 N35790 0 diode
R35791 N35790 N35791 10
D35791 N35791 0 diode
R35792 N35791 N35792 10
D35792 N35792 0 diode
R35793 N35792 N35793 10
D35793 N35793 0 diode
R35794 N35793 N35794 10
D35794 N35794 0 diode
R35795 N35794 N35795 10
D35795 N35795 0 diode
R35796 N35795 N35796 10
D35796 N35796 0 diode
R35797 N35796 N35797 10
D35797 N35797 0 diode
R35798 N35797 N35798 10
D35798 N35798 0 diode
R35799 N35798 N35799 10
D35799 N35799 0 diode
R35800 N35799 N35800 10
D35800 N35800 0 diode
R35801 N35800 N35801 10
D35801 N35801 0 diode
R35802 N35801 N35802 10
D35802 N35802 0 diode
R35803 N35802 N35803 10
D35803 N35803 0 diode
R35804 N35803 N35804 10
D35804 N35804 0 diode
R35805 N35804 N35805 10
D35805 N35805 0 diode
R35806 N35805 N35806 10
D35806 N35806 0 diode
R35807 N35806 N35807 10
D35807 N35807 0 diode
R35808 N35807 N35808 10
D35808 N35808 0 diode
R35809 N35808 N35809 10
D35809 N35809 0 diode
R35810 N35809 N35810 10
D35810 N35810 0 diode
R35811 N35810 N35811 10
D35811 N35811 0 diode
R35812 N35811 N35812 10
D35812 N35812 0 diode
R35813 N35812 N35813 10
D35813 N35813 0 diode
R35814 N35813 N35814 10
D35814 N35814 0 diode
R35815 N35814 N35815 10
D35815 N35815 0 diode
R35816 N35815 N35816 10
D35816 N35816 0 diode
R35817 N35816 N35817 10
D35817 N35817 0 diode
R35818 N35817 N35818 10
D35818 N35818 0 diode
R35819 N35818 N35819 10
D35819 N35819 0 diode
R35820 N35819 N35820 10
D35820 N35820 0 diode
R35821 N35820 N35821 10
D35821 N35821 0 diode
R35822 N35821 N35822 10
D35822 N35822 0 diode
R35823 N35822 N35823 10
D35823 N35823 0 diode
R35824 N35823 N35824 10
D35824 N35824 0 diode
R35825 N35824 N35825 10
D35825 N35825 0 diode
R35826 N35825 N35826 10
D35826 N35826 0 diode
R35827 N35826 N35827 10
D35827 N35827 0 diode
R35828 N35827 N35828 10
D35828 N35828 0 diode
R35829 N35828 N35829 10
D35829 N35829 0 diode
R35830 N35829 N35830 10
D35830 N35830 0 diode
R35831 N35830 N35831 10
D35831 N35831 0 diode
R35832 N35831 N35832 10
D35832 N35832 0 diode
R35833 N35832 N35833 10
D35833 N35833 0 diode
R35834 N35833 N35834 10
D35834 N35834 0 diode
R35835 N35834 N35835 10
D35835 N35835 0 diode
R35836 N35835 N35836 10
D35836 N35836 0 diode
R35837 N35836 N35837 10
D35837 N35837 0 diode
R35838 N35837 N35838 10
D35838 N35838 0 diode
R35839 N35838 N35839 10
D35839 N35839 0 diode
R35840 N35839 N35840 10
D35840 N35840 0 diode
R35841 N35840 N35841 10
D35841 N35841 0 diode
R35842 N35841 N35842 10
D35842 N35842 0 diode
R35843 N35842 N35843 10
D35843 N35843 0 diode
R35844 N35843 N35844 10
D35844 N35844 0 diode
R35845 N35844 N35845 10
D35845 N35845 0 diode
R35846 N35845 N35846 10
D35846 N35846 0 diode
R35847 N35846 N35847 10
D35847 N35847 0 diode
R35848 N35847 N35848 10
D35848 N35848 0 diode
R35849 N35848 N35849 10
D35849 N35849 0 diode
R35850 N35849 N35850 10
D35850 N35850 0 diode
R35851 N35850 N35851 10
D35851 N35851 0 diode
R35852 N35851 N35852 10
D35852 N35852 0 diode
R35853 N35852 N35853 10
D35853 N35853 0 diode
R35854 N35853 N35854 10
D35854 N35854 0 diode
R35855 N35854 N35855 10
D35855 N35855 0 diode
R35856 N35855 N35856 10
D35856 N35856 0 diode
R35857 N35856 N35857 10
D35857 N35857 0 diode
R35858 N35857 N35858 10
D35858 N35858 0 diode
R35859 N35858 N35859 10
D35859 N35859 0 diode
R35860 N35859 N35860 10
D35860 N35860 0 diode
R35861 N35860 N35861 10
D35861 N35861 0 diode
R35862 N35861 N35862 10
D35862 N35862 0 diode
R35863 N35862 N35863 10
D35863 N35863 0 diode
R35864 N35863 N35864 10
D35864 N35864 0 diode
R35865 N35864 N35865 10
D35865 N35865 0 diode
R35866 N35865 N35866 10
D35866 N35866 0 diode
R35867 N35866 N35867 10
D35867 N35867 0 diode
R35868 N35867 N35868 10
D35868 N35868 0 diode
R35869 N35868 N35869 10
D35869 N35869 0 diode
R35870 N35869 N35870 10
D35870 N35870 0 diode
R35871 N35870 N35871 10
D35871 N35871 0 diode
R35872 N35871 N35872 10
D35872 N35872 0 diode
R35873 N35872 N35873 10
D35873 N35873 0 diode
R35874 N35873 N35874 10
D35874 N35874 0 diode
R35875 N35874 N35875 10
D35875 N35875 0 diode
R35876 N35875 N35876 10
D35876 N35876 0 diode
R35877 N35876 N35877 10
D35877 N35877 0 diode
R35878 N35877 N35878 10
D35878 N35878 0 diode
R35879 N35878 N35879 10
D35879 N35879 0 diode
R35880 N35879 N35880 10
D35880 N35880 0 diode
R35881 N35880 N35881 10
D35881 N35881 0 diode
R35882 N35881 N35882 10
D35882 N35882 0 diode
R35883 N35882 N35883 10
D35883 N35883 0 diode
R35884 N35883 N35884 10
D35884 N35884 0 diode
R35885 N35884 N35885 10
D35885 N35885 0 diode
R35886 N35885 N35886 10
D35886 N35886 0 diode
R35887 N35886 N35887 10
D35887 N35887 0 diode
R35888 N35887 N35888 10
D35888 N35888 0 diode
R35889 N35888 N35889 10
D35889 N35889 0 diode
R35890 N35889 N35890 10
D35890 N35890 0 diode
R35891 N35890 N35891 10
D35891 N35891 0 diode
R35892 N35891 N35892 10
D35892 N35892 0 diode
R35893 N35892 N35893 10
D35893 N35893 0 diode
R35894 N35893 N35894 10
D35894 N35894 0 diode
R35895 N35894 N35895 10
D35895 N35895 0 diode
R35896 N35895 N35896 10
D35896 N35896 0 diode
R35897 N35896 N35897 10
D35897 N35897 0 diode
R35898 N35897 N35898 10
D35898 N35898 0 diode
R35899 N35898 N35899 10
D35899 N35899 0 diode
R35900 N35899 N35900 10
D35900 N35900 0 diode
R35901 N35900 N35901 10
D35901 N35901 0 diode
R35902 N35901 N35902 10
D35902 N35902 0 diode
R35903 N35902 N35903 10
D35903 N35903 0 diode
R35904 N35903 N35904 10
D35904 N35904 0 diode
R35905 N35904 N35905 10
D35905 N35905 0 diode
R35906 N35905 N35906 10
D35906 N35906 0 diode
R35907 N35906 N35907 10
D35907 N35907 0 diode
R35908 N35907 N35908 10
D35908 N35908 0 diode
R35909 N35908 N35909 10
D35909 N35909 0 diode
R35910 N35909 N35910 10
D35910 N35910 0 diode
R35911 N35910 N35911 10
D35911 N35911 0 diode
R35912 N35911 N35912 10
D35912 N35912 0 diode
R35913 N35912 N35913 10
D35913 N35913 0 diode
R35914 N35913 N35914 10
D35914 N35914 0 diode
R35915 N35914 N35915 10
D35915 N35915 0 diode
R35916 N35915 N35916 10
D35916 N35916 0 diode
R35917 N35916 N35917 10
D35917 N35917 0 diode
R35918 N35917 N35918 10
D35918 N35918 0 diode
R35919 N35918 N35919 10
D35919 N35919 0 diode
R35920 N35919 N35920 10
D35920 N35920 0 diode
R35921 N35920 N35921 10
D35921 N35921 0 diode
R35922 N35921 N35922 10
D35922 N35922 0 diode
R35923 N35922 N35923 10
D35923 N35923 0 diode
R35924 N35923 N35924 10
D35924 N35924 0 diode
R35925 N35924 N35925 10
D35925 N35925 0 diode
R35926 N35925 N35926 10
D35926 N35926 0 diode
R35927 N35926 N35927 10
D35927 N35927 0 diode
R35928 N35927 N35928 10
D35928 N35928 0 diode
R35929 N35928 N35929 10
D35929 N35929 0 diode
R35930 N35929 N35930 10
D35930 N35930 0 diode
R35931 N35930 N35931 10
D35931 N35931 0 diode
R35932 N35931 N35932 10
D35932 N35932 0 diode
R35933 N35932 N35933 10
D35933 N35933 0 diode
R35934 N35933 N35934 10
D35934 N35934 0 diode
R35935 N35934 N35935 10
D35935 N35935 0 diode
R35936 N35935 N35936 10
D35936 N35936 0 diode
R35937 N35936 N35937 10
D35937 N35937 0 diode
R35938 N35937 N35938 10
D35938 N35938 0 diode
R35939 N35938 N35939 10
D35939 N35939 0 diode
R35940 N35939 N35940 10
D35940 N35940 0 diode
R35941 N35940 N35941 10
D35941 N35941 0 diode
R35942 N35941 N35942 10
D35942 N35942 0 diode
R35943 N35942 N35943 10
D35943 N35943 0 diode
R35944 N35943 N35944 10
D35944 N35944 0 diode
R35945 N35944 N35945 10
D35945 N35945 0 diode
R35946 N35945 N35946 10
D35946 N35946 0 diode
R35947 N35946 N35947 10
D35947 N35947 0 diode
R35948 N35947 N35948 10
D35948 N35948 0 diode
R35949 N35948 N35949 10
D35949 N35949 0 diode
R35950 N35949 N35950 10
D35950 N35950 0 diode
R35951 N35950 N35951 10
D35951 N35951 0 diode
R35952 N35951 N35952 10
D35952 N35952 0 diode
R35953 N35952 N35953 10
D35953 N35953 0 diode
R35954 N35953 N35954 10
D35954 N35954 0 diode
R35955 N35954 N35955 10
D35955 N35955 0 diode
R35956 N35955 N35956 10
D35956 N35956 0 diode
R35957 N35956 N35957 10
D35957 N35957 0 diode
R35958 N35957 N35958 10
D35958 N35958 0 diode
R35959 N35958 N35959 10
D35959 N35959 0 diode
R35960 N35959 N35960 10
D35960 N35960 0 diode
R35961 N35960 N35961 10
D35961 N35961 0 diode
R35962 N35961 N35962 10
D35962 N35962 0 diode
R35963 N35962 N35963 10
D35963 N35963 0 diode
R35964 N35963 N35964 10
D35964 N35964 0 diode
R35965 N35964 N35965 10
D35965 N35965 0 diode
R35966 N35965 N35966 10
D35966 N35966 0 diode
R35967 N35966 N35967 10
D35967 N35967 0 diode
R35968 N35967 N35968 10
D35968 N35968 0 diode
R35969 N35968 N35969 10
D35969 N35969 0 diode
R35970 N35969 N35970 10
D35970 N35970 0 diode
R35971 N35970 N35971 10
D35971 N35971 0 diode
R35972 N35971 N35972 10
D35972 N35972 0 diode
R35973 N35972 N35973 10
D35973 N35973 0 diode
R35974 N35973 N35974 10
D35974 N35974 0 diode
R35975 N35974 N35975 10
D35975 N35975 0 diode
R35976 N35975 N35976 10
D35976 N35976 0 diode
R35977 N35976 N35977 10
D35977 N35977 0 diode
R35978 N35977 N35978 10
D35978 N35978 0 diode
R35979 N35978 N35979 10
D35979 N35979 0 diode
R35980 N35979 N35980 10
D35980 N35980 0 diode
R35981 N35980 N35981 10
D35981 N35981 0 diode
R35982 N35981 N35982 10
D35982 N35982 0 diode
R35983 N35982 N35983 10
D35983 N35983 0 diode
R35984 N35983 N35984 10
D35984 N35984 0 diode
R35985 N35984 N35985 10
D35985 N35985 0 diode
R35986 N35985 N35986 10
D35986 N35986 0 diode
R35987 N35986 N35987 10
D35987 N35987 0 diode
R35988 N35987 N35988 10
D35988 N35988 0 diode
R35989 N35988 N35989 10
D35989 N35989 0 diode
R35990 N35989 N35990 10
D35990 N35990 0 diode
R35991 N35990 N35991 10
D35991 N35991 0 diode
R35992 N35991 N35992 10
D35992 N35992 0 diode
R35993 N35992 N35993 10
D35993 N35993 0 diode
R35994 N35993 N35994 10
D35994 N35994 0 diode
R35995 N35994 N35995 10
D35995 N35995 0 diode
R35996 N35995 N35996 10
D35996 N35996 0 diode
R35997 N35996 N35997 10
D35997 N35997 0 diode
R35998 N35997 N35998 10
D35998 N35998 0 diode
R35999 N35998 N35999 10
D35999 N35999 0 diode
R36000 N35999 N36000 10
D36000 N36000 0 diode
R36001 N36000 N36001 10
D36001 N36001 0 diode
R36002 N36001 N36002 10
D36002 N36002 0 diode
R36003 N36002 N36003 10
D36003 N36003 0 diode
R36004 N36003 N36004 10
D36004 N36004 0 diode
R36005 N36004 N36005 10
D36005 N36005 0 diode
R36006 N36005 N36006 10
D36006 N36006 0 diode
R36007 N36006 N36007 10
D36007 N36007 0 diode
R36008 N36007 N36008 10
D36008 N36008 0 diode
R36009 N36008 N36009 10
D36009 N36009 0 diode
R36010 N36009 N36010 10
D36010 N36010 0 diode
R36011 N36010 N36011 10
D36011 N36011 0 diode
R36012 N36011 N36012 10
D36012 N36012 0 diode
R36013 N36012 N36013 10
D36013 N36013 0 diode
R36014 N36013 N36014 10
D36014 N36014 0 diode
R36015 N36014 N36015 10
D36015 N36015 0 diode
R36016 N36015 N36016 10
D36016 N36016 0 diode
R36017 N36016 N36017 10
D36017 N36017 0 diode
R36018 N36017 N36018 10
D36018 N36018 0 diode
R36019 N36018 N36019 10
D36019 N36019 0 diode
R36020 N36019 N36020 10
D36020 N36020 0 diode
R36021 N36020 N36021 10
D36021 N36021 0 diode
R36022 N36021 N36022 10
D36022 N36022 0 diode
R36023 N36022 N36023 10
D36023 N36023 0 diode
R36024 N36023 N36024 10
D36024 N36024 0 diode
R36025 N36024 N36025 10
D36025 N36025 0 diode
R36026 N36025 N36026 10
D36026 N36026 0 diode
R36027 N36026 N36027 10
D36027 N36027 0 diode
R36028 N36027 N36028 10
D36028 N36028 0 diode
R36029 N36028 N36029 10
D36029 N36029 0 diode
R36030 N36029 N36030 10
D36030 N36030 0 diode
R36031 N36030 N36031 10
D36031 N36031 0 diode
R36032 N36031 N36032 10
D36032 N36032 0 diode
R36033 N36032 N36033 10
D36033 N36033 0 diode
R36034 N36033 N36034 10
D36034 N36034 0 diode
R36035 N36034 N36035 10
D36035 N36035 0 diode
R36036 N36035 N36036 10
D36036 N36036 0 diode
R36037 N36036 N36037 10
D36037 N36037 0 diode
R36038 N36037 N36038 10
D36038 N36038 0 diode
R36039 N36038 N36039 10
D36039 N36039 0 diode
R36040 N36039 N36040 10
D36040 N36040 0 diode
R36041 N36040 N36041 10
D36041 N36041 0 diode
R36042 N36041 N36042 10
D36042 N36042 0 diode
R36043 N36042 N36043 10
D36043 N36043 0 diode
R36044 N36043 N36044 10
D36044 N36044 0 diode
R36045 N36044 N36045 10
D36045 N36045 0 diode
R36046 N36045 N36046 10
D36046 N36046 0 diode
R36047 N36046 N36047 10
D36047 N36047 0 diode
R36048 N36047 N36048 10
D36048 N36048 0 diode
R36049 N36048 N36049 10
D36049 N36049 0 diode
R36050 N36049 N36050 10
D36050 N36050 0 diode
R36051 N36050 N36051 10
D36051 N36051 0 diode
R36052 N36051 N36052 10
D36052 N36052 0 diode
R36053 N36052 N36053 10
D36053 N36053 0 diode
R36054 N36053 N36054 10
D36054 N36054 0 diode
R36055 N36054 N36055 10
D36055 N36055 0 diode
R36056 N36055 N36056 10
D36056 N36056 0 diode
R36057 N36056 N36057 10
D36057 N36057 0 diode
R36058 N36057 N36058 10
D36058 N36058 0 diode
R36059 N36058 N36059 10
D36059 N36059 0 diode
R36060 N36059 N36060 10
D36060 N36060 0 diode
R36061 N36060 N36061 10
D36061 N36061 0 diode
R36062 N36061 N36062 10
D36062 N36062 0 diode
R36063 N36062 N36063 10
D36063 N36063 0 diode
R36064 N36063 N36064 10
D36064 N36064 0 diode
R36065 N36064 N36065 10
D36065 N36065 0 diode
R36066 N36065 N36066 10
D36066 N36066 0 diode
R36067 N36066 N36067 10
D36067 N36067 0 diode
R36068 N36067 N36068 10
D36068 N36068 0 diode
R36069 N36068 N36069 10
D36069 N36069 0 diode
R36070 N36069 N36070 10
D36070 N36070 0 diode
R36071 N36070 N36071 10
D36071 N36071 0 diode
R36072 N36071 N36072 10
D36072 N36072 0 diode
R36073 N36072 N36073 10
D36073 N36073 0 diode
R36074 N36073 N36074 10
D36074 N36074 0 diode
R36075 N36074 N36075 10
D36075 N36075 0 diode
R36076 N36075 N36076 10
D36076 N36076 0 diode
R36077 N36076 N36077 10
D36077 N36077 0 diode
R36078 N36077 N36078 10
D36078 N36078 0 diode
R36079 N36078 N36079 10
D36079 N36079 0 diode
R36080 N36079 N36080 10
D36080 N36080 0 diode
R36081 N36080 N36081 10
D36081 N36081 0 diode
R36082 N36081 N36082 10
D36082 N36082 0 diode
R36083 N36082 N36083 10
D36083 N36083 0 diode
R36084 N36083 N36084 10
D36084 N36084 0 diode
R36085 N36084 N36085 10
D36085 N36085 0 diode
R36086 N36085 N36086 10
D36086 N36086 0 diode
R36087 N36086 N36087 10
D36087 N36087 0 diode
R36088 N36087 N36088 10
D36088 N36088 0 diode
R36089 N36088 N36089 10
D36089 N36089 0 diode
R36090 N36089 N36090 10
D36090 N36090 0 diode
R36091 N36090 N36091 10
D36091 N36091 0 diode
R36092 N36091 N36092 10
D36092 N36092 0 diode
R36093 N36092 N36093 10
D36093 N36093 0 diode
R36094 N36093 N36094 10
D36094 N36094 0 diode
R36095 N36094 N36095 10
D36095 N36095 0 diode
R36096 N36095 N36096 10
D36096 N36096 0 diode
R36097 N36096 N36097 10
D36097 N36097 0 diode
R36098 N36097 N36098 10
D36098 N36098 0 diode
R36099 N36098 N36099 10
D36099 N36099 0 diode
R36100 N36099 N36100 10
D36100 N36100 0 diode
R36101 N36100 N36101 10
D36101 N36101 0 diode
R36102 N36101 N36102 10
D36102 N36102 0 diode
R36103 N36102 N36103 10
D36103 N36103 0 diode
R36104 N36103 N36104 10
D36104 N36104 0 diode
R36105 N36104 N36105 10
D36105 N36105 0 diode
R36106 N36105 N36106 10
D36106 N36106 0 diode
R36107 N36106 N36107 10
D36107 N36107 0 diode
R36108 N36107 N36108 10
D36108 N36108 0 diode
R36109 N36108 N36109 10
D36109 N36109 0 diode
R36110 N36109 N36110 10
D36110 N36110 0 diode
R36111 N36110 N36111 10
D36111 N36111 0 diode
R36112 N36111 N36112 10
D36112 N36112 0 diode
R36113 N36112 N36113 10
D36113 N36113 0 diode
R36114 N36113 N36114 10
D36114 N36114 0 diode
R36115 N36114 N36115 10
D36115 N36115 0 diode
R36116 N36115 N36116 10
D36116 N36116 0 diode
R36117 N36116 N36117 10
D36117 N36117 0 diode
R36118 N36117 N36118 10
D36118 N36118 0 diode
R36119 N36118 N36119 10
D36119 N36119 0 diode
R36120 N36119 N36120 10
D36120 N36120 0 diode
R36121 N36120 N36121 10
D36121 N36121 0 diode
R36122 N36121 N36122 10
D36122 N36122 0 diode
R36123 N36122 N36123 10
D36123 N36123 0 diode
R36124 N36123 N36124 10
D36124 N36124 0 diode
R36125 N36124 N36125 10
D36125 N36125 0 diode
R36126 N36125 N36126 10
D36126 N36126 0 diode
R36127 N36126 N36127 10
D36127 N36127 0 diode
R36128 N36127 N36128 10
D36128 N36128 0 diode
R36129 N36128 N36129 10
D36129 N36129 0 diode
R36130 N36129 N36130 10
D36130 N36130 0 diode
R36131 N36130 N36131 10
D36131 N36131 0 diode
R36132 N36131 N36132 10
D36132 N36132 0 diode
R36133 N36132 N36133 10
D36133 N36133 0 diode
R36134 N36133 N36134 10
D36134 N36134 0 diode
R36135 N36134 N36135 10
D36135 N36135 0 diode
R36136 N36135 N36136 10
D36136 N36136 0 diode
R36137 N36136 N36137 10
D36137 N36137 0 diode
R36138 N36137 N36138 10
D36138 N36138 0 diode
R36139 N36138 N36139 10
D36139 N36139 0 diode
R36140 N36139 N36140 10
D36140 N36140 0 diode
R36141 N36140 N36141 10
D36141 N36141 0 diode
R36142 N36141 N36142 10
D36142 N36142 0 diode
R36143 N36142 N36143 10
D36143 N36143 0 diode
R36144 N36143 N36144 10
D36144 N36144 0 diode
R36145 N36144 N36145 10
D36145 N36145 0 diode
R36146 N36145 N36146 10
D36146 N36146 0 diode
R36147 N36146 N36147 10
D36147 N36147 0 diode
R36148 N36147 N36148 10
D36148 N36148 0 diode
R36149 N36148 N36149 10
D36149 N36149 0 diode
R36150 N36149 N36150 10
D36150 N36150 0 diode
R36151 N36150 N36151 10
D36151 N36151 0 diode
R36152 N36151 N36152 10
D36152 N36152 0 diode
R36153 N36152 N36153 10
D36153 N36153 0 diode
R36154 N36153 N36154 10
D36154 N36154 0 diode
R36155 N36154 N36155 10
D36155 N36155 0 diode
R36156 N36155 N36156 10
D36156 N36156 0 diode
R36157 N36156 N36157 10
D36157 N36157 0 diode
R36158 N36157 N36158 10
D36158 N36158 0 diode
R36159 N36158 N36159 10
D36159 N36159 0 diode
R36160 N36159 N36160 10
D36160 N36160 0 diode
R36161 N36160 N36161 10
D36161 N36161 0 diode
R36162 N36161 N36162 10
D36162 N36162 0 diode
R36163 N36162 N36163 10
D36163 N36163 0 diode
R36164 N36163 N36164 10
D36164 N36164 0 diode
R36165 N36164 N36165 10
D36165 N36165 0 diode
R36166 N36165 N36166 10
D36166 N36166 0 diode
R36167 N36166 N36167 10
D36167 N36167 0 diode
R36168 N36167 N36168 10
D36168 N36168 0 diode
R36169 N36168 N36169 10
D36169 N36169 0 diode
R36170 N36169 N36170 10
D36170 N36170 0 diode
R36171 N36170 N36171 10
D36171 N36171 0 diode
R36172 N36171 N36172 10
D36172 N36172 0 diode
R36173 N36172 N36173 10
D36173 N36173 0 diode
R36174 N36173 N36174 10
D36174 N36174 0 diode
R36175 N36174 N36175 10
D36175 N36175 0 diode
R36176 N36175 N36176 10
D36176 N36176 0 diode
R36177 N36176 N36177 10
D36177 N36177 0 diode
R36178 N36177 N36178 10
D36178 N36178 0 diode
R36179 N36178 N36179 10
D36179 N36179 0 diode
R36180 N36179 N36180 10
D36180 N36180 0 diode
R36181 N36180 N36181 10
D36181 N36181 0 diode
R36182 N36181 N36182 10
D36182 N36182 0 diode
R36183 N36182 N36183 10
D36183 N36183 0 diode
R36184 N36183 N36184 10
D36184 N36184 0 diode
R36185 N36184 N36185 10
D36185 N36185 0 diode
R36186 N36185 N36186 10
D36186 N36186 0 diode
R36187 N36186 N36187 10
D36187 N36187 0 diode
R36188 N36187 N36188 10
D36188 N36188 0 diode
R36189 N36188 N36189 10
D36189 N36189 0 diode
R36190 N36189 N36190 10
D36190 N36190 0 diode
R36191 N36190 N36191 10
D36191 N36191 0 diode
R36192 N36191 N36192 10
D36192 N36192 0 diode
R36193 N36192 N36193 10
D36193 N36193 0 diode
R36194 N36193 N36194 10
D36194 N36194 0 diode
R36195 N36194 N36195 10
D36195 N36195 0 diode
R36196 N36195 N36196 10
D36196 N36196 0 diode
R36197 N36196 N36197 10
D36197 N36197 0 diode
R36198 N36197 N36198 10
D36198 N36198 0 diode
R36199 N36198 N36199 10
D36199 N36199 0 diode
R36200 N36199 N36200 10
D36200 N36200 0 diode
R36201 N36200 N36201 10
D36201 N36201 0 diode
R36202 N36201 N36202 10
D36202 N36202 0 diode
R36203 N36202 N36203 10
D36203 N36203 0 diode
R36204 N36203 N36204 10
D36204 N36204 0 diode
R36205 N36204 N36205 10
D36205 N36205 0 diode
R36206 N36205 N36206 10
D36206 N36206 0 diode
R36207 N36206 N36207 10
D36207 N36207 0 diode
R36208 N36207 N36208 10
D36208 N36208 0 diode
R36209 N36208 N36209 10
D36209 N36209 0 diode
R36210 N36209 N36210 10
D36210 N36210 0 diode
R36211 N36210 N36211 10
D36211 N36211 0 diode
R36212 N36211 N36212 10
D36212 N36212 0 diode
R36213 N36212 N36213 10
D36213 N36213 0 diode
R36214 N36213 N36214 10
D36214 N36214 0 diode
R36215 N36214 N36215 10
D36215 N36215 0 diode
R36216 N36215 N36216 10
D36216 N36216 0 diode
R36217 N36216 N36217 10
D36217 N36217 0 diode
R36218 N36217 N36218 10
D36218 N36218 0 diode
R36219 N36218 N36219 10
D36219 N36219 0 diode
R36220 N36219 N36220 10
D36220 N36220 0 diode
R36221 N36220 N36221 10
D36221 N36221 0 diode
R36222 N36221 N36222 10
D36222 N36222 0 diode
R36223 N36222 N36223 10
D36223 N36223 0 diode
R36224 N36223 N36224 10
D36224 N36224 0 diode
R36225 N36224 N36225 10
D36225 N36225 0 diode
R36226 N36225 N36226 10
D36226 N36226 0 diode
R36227 N36226 N36227 10
D36227 N36227 0 diode
R36228 N36227 N36228 10
D36228 N36228 0 diode
R36229 N36228 N36229 10
D36229 N36229 0 diode
R36230 N36229 N36230 10
D36230 N36230 0 diode
R36231 N36230 N36231 10
D36231 N36231 0 diode
R36232 N36231 N36232 10
D36232 N36232 0 diode
R36233 N36232 N36233 10
D36233 N36233 0 diode
R36234 N36233 N36234 10
D36234 N36234 0 diode
R36235 N36234 N36235 10
D36235 N36235 0 diode
R36236 N36235 N36236 10
D36236 N36236 0 diode
R36237 N36236 N36237 10
D36237 N36237 0 diode
R36238 N36237 N36238 10
D36238 N36238 0 diode
R36239 N36238 N36239 10
D36239 N36239 0 diode
R36240 N36239 N36240 10
D36240 N36240 0 diode
R36241 N36240 N36241 10
D36241 N36241 0 diode
R36242 N36241 N36242 10
D36242 N36242 0 diode
R36243 N36242 N36243 10
D36243 N36243 0 diode
R36244 N36243 N36244 10
D36244 N36244 0 diode
R36245 N36244 N36245 10
D36245 N36245 0 diode
R36246 N36245 N36246 10
D36246 N36246 0 diode
R36247 N36246 N36247 10
D36247 N36247 0 diode
R36248 N36247 N36248 10
D36248 N36248 0 diode
R36249 N36248 N36249 10
D36249 N36249 0 diode
R36250 N36249 N36250 10
D36250 N36250 0 diode
R36251 N36250 N36251 10
D36251 N36251 0 diode
R36252 N36251 N36252 10
D36252 N36252 0 diode
R36253 N36252 N36253 10
D36253 N36253 0 diode
R36254 N36253 N36254 10
D36254 N36254 0 diode
R36255 N36254 N36255 10
D36255 N36255 0 diode
R36256 N36255 N36256 10
D36256 N36256 0 diode
R36257 N36256 N36257 10
D36257 N36257 0 diode
R36258 N36257 N36258 10
D36258 N36258 0 diode
R36259 N36258 N36259 10
D36259 N36259 0 diode
R36260 N36259 N36260 10
D36260 N36260 0 diode
R36261 N36260 N36261 10
D36261 N36261 0 diode
R36262 N36261 N36262 10
D36262 N36262 0 diode
R36263 N36262 N36263 10
D36263 N36263 0 diode
R36264 N36263 N36264 10
D36264 N36264 0 diode
R36265 N36264 N36265 10
D36265 N36265 0 diode
R36266 N36265 N36266 10
D36266 N36266 0 diode
R36267 N36266 N36267 10
D36267 N36267 0 diode
R36268 N36267 N36268 10
D36268 N36268 0 diode
R36269 N36268 N36269 10
D36269 N36269 0 diode
R36270 N36269 N36270 10
D36270 N36270 0 diode
R36271 N36270 N36271 10
D36271 N36271 0 diode
R36272 N36271 N36272 10
D36272 N36272 0 diode
R36273 N36272 N36273 10
D36273 N36273 0 diode
R36274 N36273 N36274 10
D36274 N36274 0 diode
R36275 N36274 N36275 10
D36275 N36275 0 diode
R36276 N36275 N36276 10
D36276 N36276 0 diode
R36277 N36276 N36277 10
D36277 N36277 0 diode
R36278 N36277 N36278 10
D36278 N36278 0 diode
R36279 N36278 N36279 10
D36279 N36279 0 diode
R36280 N36279 N36280 10
D36280 N36280 0 diode
R36281 N36280 N36281 10
D36281 N36281 0 diode
R36282 N36281 N36282 10
D36282 N36282 0 diode
R36283 N36282 N36283 10
D36283 N36283 0 diode
R36284 N36283 N36284 10
D36284 N36284 0 diode
R36285 N36284 N36285 10
D36285 N36285 0 diode
R36286 N36285 N36286 10
D36286 N36286 0 diode
R36287 N36286 N36287 10
D36287 N36287 0 diode
R36288 N36287 N36288 10
D36288 N36288 0 diode
R36289 N36288 N36289 10
D36289 N36289 0 diode
R36290 N36289 N36290 10
D36290 N36290 0 diode
R36291 N36290 N36291 10
D36291 N36291 0 diode
R36292 N36291 N36292 10
D36292 N36292 0 diode
R36293 N36292 N36293 10
D36293 N36293 0 diode
R36294 N36293 N36294 10
D36294 N36294 0 diode
R36295 N36294 N36295 10
D36295 N36295 0 diode
R36296 N36295 N36296 10
D36296 N36296 0 diode
R36297 N36296 N36297 10
D36297 N36297 0 diode
R36298 N36297 N36298 10
D36298 N36298 0 diode
R36299 N36298 N36299 10
D36299 N36299 0 diode
R36300 N36299 N36300 10
D36300 N36300 0 diode
R36301 N36300 N36301 10
D36301 N36301 0 diode
R36302 N36301 N36302 10
D36302 N36302 0 diode
R36303 N36302 N36303 10
D36303 N36303 0 diode
R36304 N36303 N36304 10
D36304 N36304 0 diode
R36305 N36304 N36305 10
D36305 N36305 0 diode
R36306 N36305 N36306 10
D36306 N36306 0 diode
R36307 N36306 N36307 10
D36307 N36307 0 diode
R36308 N36307 N36308 10
D36308 N36308 0 diode
R36309 N36308 N36309 10
D36309 N36309 0 diode
R36310 N36309 N36310 10
D36310 N36310 0 diode
R36311 N36310 N36311 10
D36311 N36311 0 diode
R36312 N36311 N36312 10
D36312 N36312 0 diode
R36313 N36312 N36313 10
D36313 N36313 0 diode
R36314 N36313 N36314 10
D36314 N36314 0 diode
R36315 N36314 N36315 10
D36315 N36315 0 diode
R36316 N36315 N36316 10
D36316 N36316 0 diode
R36317 N36316 N36317 10
D36317 N36317 0 diode
R36318 N36317 N36318 10
D36318 N36318 0 diode
R36319 N36318 N36319 10
D36319 N36319 0 diode
R36320 N36319 N36320 10
D36320 N36320 0 diode
R36321 N36320 N36321 10
D36321 N36321 0 diode
R36322 N36321 N36322 10
D36322 N36322 0 diode
R36323 N36322 N36323 10
D36323 N36323 0 diode
R36324 N36323 N36324 10
D36324 N36324 0 diode
R36325 N36324 N36325 10
D36325 N36325 0 diode
R36326 N36325 N36326 10
D36326 N36326 0 diode
R36327 N36326 N36327 10
D36327 N36327 0 diode
R36328 N36327 N36328 10
D36328 N36328 0 diode
R36329 N36328 N36329 10
D36329 N36329 0 diode
R36330 N36329 N36330 10
D36330 N36330 0 diode
R36331 N36330 N36331 10
D36331 N36331 0 diode
R36332 N36331 N36332 10
D36332 N36332 0 diode
R36333 N36332 N36333 10
D36333 N36333 0 diode
R36334 N36333 N36334 10
D36334 N36334 0 diode
R36335 N36334 N36335 10
D36335 N36335 0 diode
R36336 N36335 N36336 10
D36336 N36336 0 diode
R36337 N36336 N36337 10
D36337 N36337 0 diode
R36338 N36337 N36338 10
D36338 N36338 0 diode
R36339 N36338 N36339 10
D36339 N36339 0 diode
R36340 N36339 N36340 10
D36340 N36340 0 diode
R36341 N36340 N36341 10
D36341 N36341 0 diode
R36342 N36341 N36342 10
D36342 N36342 0 diode
R36343 N36342 N36343 10
D36343 N36343 0 diode
R36344 N36343 N36344 10
D36344 N36344 0 diode
R36345 N36344 N36345 10
D36345 N36345 0 diode
R36346 N36345 N36346 10
D36346 N36346 0 diode
R36347 N36346 N36347 10
D36347 N36347 0 diode
R36348 N36347 N36348 10
D36348 N36348 0 diode
R36349 N36348 N36349 10
D36349 N36349 0 diode
R36350 N36349 N36350 10
D36350 N36350 0 diode
R36351 N36350 N36351 10
D36351 N36351 0 diode
R36352 N36351 N36352 10
D36352 N36352 0 diode
R36353 N36352 N36353 10
D36353 N36353 0 diode
R36354 N36353 N36354 10
D36354 N36354 0 diode
R36355 N36354 N36355 10
D36355 N36355 0 diode
R36356 N36355 N36356 10
D36356 N36356 0 diode
R36357 N36356 N36357 10
D36357 N36357 0 diode
R36358 N36357 N36358 10
D36358 N36358 0 diode
R36359 N36358 N36359 10
D36359 N36359 0 diode
R36360 N36359 N36360 10
D36360 N36360 0 diode
R36361 N36360 N36361 10
D36361 N36361 0 diode
R36362 N36361 N36362 10
D36362 N36362 0 diode
R36363 N36362 N36363 10
D36363 N36363 0 diode
R36364 N36363 N36364 10
D36364 N36364 0 diode
R36365 N36364 N36365 10
D36365 N36365 0 diode
R36366 N36365 N36366 10
D36366 N36366 0 diode
R36367 N36366 N36367 10
D36367 N36367 0 diode
R36368 N36367 N36368 10
D36368 N36368 0 diode
R36369 N36368 N36369 10
D36369 N36369 0 diode
R36370 N36369 N36370 10
D36370 N36370 0 diode
R36371 N36370 N36371 10
D36371 N36371 0 diode
R36372 N36371 N36372 10
D36372 N36372 0 diode
R36373 N36372 N36373 10
D36373 N36373 0 diode
R36374 N36373 N36374 10
D36374 N36374 0 diode
R36375 N36374 N36375 10
D36375 N36375 0 diode
R36376 N36375 N36376 10
D36376 N36376 0 diode
R36377 N36376 N36377 10
D36377 N36377 0 diode
R36378 N36377 N36378 10
D36378 N36378 0 diode
R36379 N36378 N36379 10
D36379 N36379 0 diode
R36380 N36379 N36380 10
D36380 N36380 0 diode
R36381 N36380 N36381 10
D36381 N36381 0 diode
R36382 N36381 N36382 10
D36382 N36382 0 diode
R36383 N36382 N36383 10
D36383 N36383 0 diode
R36384 N36383 N36384 10
D36384 N36384 0 diode
R36385 N36384 N36385 10
D36385 N36385 0 diode
R36386 N36385 N36386 10
D36386 N36386 0 diode
R36387 N36386 N36387 10
D36387 N36387 0 diode
R36388 N36387 N36388 10
D36388 N36388 0 diode
R36389 N36388 N36389 10
D36389 N36389 0 diode
R36390 N36389 N36390 10
D36390 N36390 0 diode
R36391 N36390 N36391 10
D36391 N36391 0 diode
R36392 N36391 N36392 10
D36392 N36392 0 diode
R36393 N36392 N36393 10
D36393 N36393 0 diode
R36394 N36393 N36394 10
D36394 N36394 0 diode
R36395 N36394 N36395 10
D36395 N36395 0 diode
R36396 N36395 N36396 10
D36396 N36396 0 diode
R36397 N36396 N36397 10
D36397 N36397 0 diode
R36398 N36397 N36398 10
D36398 N36398 0 diode
R36399 N36398 N36399 10
D36399 N36399 0 diode
R36400 N36399 N36400 10
D36400 N36400 0 diode
R36401 N36400 N36401 10
D36401 N36401 0 diode
R36402 N36401 N36402 10
D36402 N36402 0 diode
R36403 N36402 N36403 10
D36403 N36403 0 diode
R36404 N36403 N36404 10
D36404 N36404 0 diode
R36405 N36404 N36405 10
D36405 N36405 0 diode
R36406 N36405 N36406 10
D36406 N36406 0 diode
R36407 N36406 N36407 10
D36407 N36407 0 diode
R36408 N36407 N36408 10
D36408 N36408 0 diode
R36409 N36408 N36409 10
D36409 N36409 0 diode
R36410 N36409 N36410 10
D36410 N36410 0 diode
R36411 N36410 N36411 10
D36411 N36411 0 diode
R36412 N36411 N36412 10
D36412 N36412 0 diode
R36413 N36412 N36413 10
D36413 N36413 0 diode
R36414 N36413 N36414 10
D36414 N36414 0 diode
R36415 N36414 N36415 10
D36415 N36415 0 diode
R36416 N36415 N36416 10
D36416 N36416 0 diode
R36417 N36416 N36417 10
D36417 N36417 0 diode
R36418 N36417 N36418 10
D36418 N36418 0 diode
R36419 N36418 N36419 10
D36419 N36419 0 diode
R36420 N36419 N36420 10
D36420 N36420 0 diode
R36421 N36420 N36421 10
D36421 N36421 0 diode
R36422 N36421 N36422 10
D36422 N36422 0 diode
R36423 N36422 N36423 10
D36423 N36423 0 diode
R36424 N36423 N36424 10
D36424 N36424 0 diode
R36425 N36424 N36425 10
D36425 N36425 0 diode
R36426 N36425 N36426 10
D36426 N36426 0 diode
R36427 N36426 N36427 10
D36427 N36427 0 diode
R36428 N36427 N36428 10
D36428 N36428 0 diode
R36429 N36428 N36429 10
D36429 N36429 0 diode
R36430 N36429 N36430 10
D36430 N36430 0 diode
R36431 N36430 N36431 10
D36431 N36431 0 diode
R36432 N36431 N36432 10
D36432 N36432 0 diode
R36433 N36432 N36433 10
D36433 N36433 0 diode
R36434 N36433 N36434 10
D36434 N36434 0 diode
R36435 N36434 N36435 10
D36435 N36435 0 diode
R36436 N36435 N36436 10
D36436 N36436 0 diode
R36437 N36436 N36437 10
D36437 N36437 0 diode
R36438 N36437 N36438 10
D36438 N36438 0 diode
R36439 N36438 N36439 10
D36439 N36439 0 diode
R36440 N36439 N36440 10
D36440 N36440 0 diode
R36441 N36440 N36441 10
D36441 N36441 0 diode
R36442 N36441 N36442 10
D36442 N36442 0 diode
R36443 N36442 N36443 10
D36443 N36443 0 diode
R36444 N36443 N36444 10
D36444 N36444 0 diode
R36445 N36444 N36445 10
D36445 N36445 0 diode
R36446 N36445 N36446 10
D36446 N36446 0 diode
R36447 N36446 N36447 10
D36447 N36447 0 diode
R36448 N36447 N36448 10
D36448 N36448 0 diode
R36449 N36448 N36449 10
D36449 N36449 0 diode
R36450 N36449 N36450 10
D36450 N36450 0 diode
R36451 N36450 N36451 10
D36451 N36451 0 diode
R36452 N36451 N36452 10
D36452 N36452 0 diode
R36453 N36452 N36453 10
D36453 N36453 0 diode
R36454 N36453 N36454 10
D36454 N36454 0 diode
R36455 N36454 N36455 10
D36455 N36455 0 diode
R36456 N36455 N36456 10
D36456 N36456 0 diode
R36457 N36456 N36457 10
D36457 N36457 0 diode
R36458 N36457 N36458 10
D36458 N36458 0 diode
R36459 N36458 N36459 10
D36459 N36459 0 diode
R36460 N36459 N36460 10
D36460 N36460 0 diode
R36461 N36460 N36461 10
D36461 N36461 0 diode
R36462 N36461 N36462 10
D36462 N36462 0 diode
R36463 N36462 N36463 10
D36463 N36463 0 diode
R36464 N36463 N36464 10
D36464 N36464 0 diode
R36465 N36464 N36465 10
D36465 N36465 0 diode
R36466 N36465 N36466 10
D36466 N36466 0 diode
R36467 N36466 N36467 10
D36467 N36467 0 diode
R36468 N36467 N36468 10
D36468 N36468 0 diode
R36469 N36468 N36469 10
D36469 N36469 0 diode
R36470 N36469 N36470 10
D36470 N36470 0 diode
R36471 N36470 N36471 10
D36471 N36471 0 diode
R36472 N36471 N36472 10
D36472 N36472 0 diode
R36473 N36472 N36473 10
D36473 N36473 0 diode
R36474 N36473 N36474 10
D36474 N36474 0 diode
R36475 N36474 N36475 10
D36475 N36475 0 diode
R36476 N36475 N36476 10
D36476 N36476 0 diode
R36477 N36476 N36477 10
D36477 N36477 0 diode
R36478 N36477 N36478 10
D36478 N36478 0 diode
R36479 N36478 N36479 10
D36479 N36479 0 diode
R36480 N36479 N36480 10
D36480 N36480 0 diode
R36481 N36480 N36481 10
D36481 N36481 0 diode
R36482 N36481 N36482 10
D36482 N36482 0 diode
R36483 N36482 N36483 10
D36483 N36483 0 diode
R36484 N36483 N36484 10
D36484 N36484 0 diode
R36485 N36484 N36485 10
D36485 N36485 0 diode
R36486 N36485 N36486 10
D36486 N36486 0 diode
R36487 N36486 N36487 10
D36487 N36487 0 diode
R36488 N36487 N36488 10
D36488 N36488 0 diode
R36489 N36488 N36489 10
D36489 N36489 0 diode
R36490 N36489 N36490 10
D36490 N36490 0 diode
R36491 N36490 N36491 10
D36491 N36491 0 diode
R36492 N36491 N36492 10
D36492 N36492 0 diode
R36493 N36492 N36493 10
D36493 N36493 0 diode
R36494 N36493 N36494 10
D36494 N36494 0 diode
R36495 N36494 N36495 10
D36495 N36495 0 diode
R36496 N36495 N36496 10
D36496 N36496 0 diode
R36497 N36496 N36497 10
D36497 N36497 0 diode
R36498 N36497 N36498 10
D36498 N36498 0 diode
R36499 N36498 N36499 10
D36499 N36499 0 diode
R36500 N36499 N36500 10
D36500 N36500 0 diode
R36501 N36500 N36501 10
D36501 N36501 0 diode
R36502 N36501 N36502 10
D36502 N36502 0 diode
R36503 N36502 N36503 10
D36503 N36503 0 diode
R36504 N36503 N36504 10
D36504 N36504 0 diode
R36505 N36504 N36505 10
D36505 N36505 0 diode
R36506 N36505 N36506 10
D36506 N36506 0 diode
R36507 N36506 N36507 10
D36507 N36507 0 diode
R36508 N36507 N36508 10
D36508 N36508 0 diode
R36509 N36508 N36509 10
D36509 N36509 0 diode
R36510 N36509 N36510 10
D36510 N36510 0 diode
R36511 N36510 N36511 10
D36511 N36511 0 diode
R36512 N36511 N36512 10
D36512 N36512 0 diode
R36513 N36512 N36513 10
D36513 N36513 0 diode
R36514 N36513 N36514 10
D36514 N36514 0 diode
R36515 N36514 N36515 10
D36515 N36515 0 diode
R36516 N36515 N36516 10
D36516 N36516 0 diode
R36517 N36516 N36517 10
D36517 N36517 0 diode
R36518 N36517 N36518 10
D36518 N36518 0 diode
R36519 N36518 N36519 10
D36519 N36519 0 diode
R36520 N36519 N36520 10
D36520 N36520 0 diode
R36521 N36520 N36521 10
D36521 N36521 0 diode
R36522 N36521 N36522 10
D36522 N36522 0 diode
R36523 N36522 N36523 10
D36523 N36523 0 diode
R36524 N36523 N36524 10
D36524 N36524 0 diode
R36525 N36524 N36525 10
D36525 N36525 0 diode
R36526 N36525 N36526 10
D36526 N36526 0 diode
R36527 N36526 N36527 10
D36527 N36527 0 diode
R36528 N36527 N36528 10
D36528 N36528 0 diode
R36529 N36528 N36529 10
D36529 N36529 0 diode
R36530 N36529 N36530 10
D36530 N36530 0 diode
R36531 N36530 N36531 10
D36531 N36531 0 diode
R36532 N36531 N36532 10
D36532 N36532 0 diode
R36533 N36532 N36533 10
D36533 N36533 0 diode
R36534 N36533 N36534 10
D36534 N36534 0 diode
R36535 N36534 N36535 10
D36535 N36535 0 diode
R36536 N36535 N36536 10
D36536 N36536 0 diode
R36537 N36536 N36537 10
D36537 N36537 0 diode
R36538 N36537 N36538 10
D36538 N36538 0 diode
R36539 N36538 N36539 10
D36539 N36539 0 diode
R36540 N36539 N36540 10
D36540 N36540 0 diode
R36541 N36540 N36541 10
D36541 N36541 0 diode
R36542 N36541 N36542 10
D36542 N36542 0 diode
R36543 N36542 N36543 10
D36543 N36543 0 diode
R36544 N36543 N36544 10
D36544 N36544 0 diode
R36545 N36544 N36545 10
D36545 N36545 0 diode
R36546 N36545 N36546 10
D36546 N36546 0 diode
R36547 N36546 N36547 10
D36547 N36547 0 diode
R36548 N36547 N36548 10
D36548 N36548 0 diode
R36549 N36548 N36549 10
D36549 N36549 0 diode
R36550 N36549 N36550 10
D36550 N36550 0 diode
R36551 N36550 N36551 10
D36551 N36551 0 diode
R36552 N36551 N36552 10
D36552 N36552 0 diode
R36553 N36552 N36553 10
D36553 N36553 0 diode
R36554 N36553 N36554 10
D36554 N36554 0 diode
R36555 N36554 N36555 10
D36555 N36555 0 diode
R36556 N36555 N36556 10
D36556 N36556 0 diode
R36557 N36556 N36557 10
D36557 N36557 0 diode
R36558 N36557 N36558 10
D36558 N36558 0 diode
R36559 N36558 N36559 10
D36559 N36559 0 diode
R36560 N36559 N36560 10
D36560 N36560 0 diode
R36561 N36560 N36561 10
D36561 N36561 0 diode
R36562 N36561 N36562 10
D36562 N36562 0 diode
R36563 N36562 N36563 10
D36563 N36563 0 diode
R36564 N36563 N36564 10
D36564 N36564 0 diode
R36565 N36564 N36565 10
D36565 N36565 0 diode
R36566 N36565 N36566 10
D36566 N36566 0 diode
R36567 N36566 N36567 10
D36567 N36567 0 diode
R36568 N36567 N36568 10
D36568 N36568 0 diode
R36569 N36568 N36569 10
D36569 N36569 0 diode
R36570 N36569 N36570 10
D36570 N36570 0 diode
R36571 N36570 N36571 10
D36571 N36571 0 diode
R36572 N36571 N36572 10
D36572 N36572 0 diode
R36573 N36572 N36573 10
D36573 N36573 0 diode
R36574 N36573 N36574 10
D36574 N36574 0 diode
R36575 N36574 N36575 10
D36575 N36575 0 diode
R36576 N36575 N36576 10
D36576 N36576 0 diode
R36577 N36576 N36577 10
D36577 N36577 0 diode
R36578 N36577 N36578 10
D36578 N36578 0 diode
R36579 N36578 N36579 10
D36579 N36579 0 diode
R36580 N36579 N36580 10
D36580 N36580 0 diode
R36581 N36580 N36581 10
D36581 N36581 0 diode
R36582 N36581 N36582 10
D36582 N36582 0 diode
R36583 N36582 N36583 10
D36583 N36583 0 diode
R36584 N36583 N36584 10
D36584 N36584 0 diode
R36585 N36584 N36585 10
D36585 N36585 0 diode
R36586 N36585 N36586 10
D36586 N36586 0 diode
R36587 N36586 N36587 10
D36587 N36587 0 diode
R36588 N36587 N36588 10
D36588 N36588 0 diode
R36589 N36588 N36589 10
D36589 N36589 0 diode
R36590 N36589 N36590 10
D36590 N36590 0 diode
R36591 N36590 N36591 10
D36591 N36591 0 diode
R36592 N36591 N36592 10
D36592 N36592 0 diode
R36593 N36592 N36593 10
D36593 N36593 0 diode
R36594 N36593 N36594 10
D36594 N36594 0 diode
R36595 N36594 N36595 10
D36595 N36595 0 diode
R36596 N36595 N36596 10
D36596 N36596 0 diode
R36597 N36596 N36597 10
D36597 N36597 0 diode
R36598 N36597 N36598 10
D36598 N36598 0 diode
R36599 N36598 N36599 10
D36599 N36599 0 diode
R36600 N36599 N36600 10
D36600 N36600 0 diode
R36601 N36600 N36601 10
D36601 N36601 0 diode
R36602 N36601 N36602 10
D36602 N36602 0 diode
R36603 N36602 N36603 10
D36603 N36603 0 diode
R36604 N36603 N36604 10
D36604 N36604 0 diode
R36605 N36604 N36605 10
D36605 N36605 0 diode
R36606 N36605 N36606 10
D36606 N36606 0 diode
R36607 N36606 N36607 10
D36607 N36607 0 diode
R36608 N36607 N36608 10
D36608 N36608 0 diode
R36609 N36608 N36609 10
D36609 N36609 0 diode
R36610 N36609 N36610 10
D36610 N36610 0 diode
R36611 N36610 N36611 10
D36611 N36611 0 diode
R36612 N36611 N36612 10
D36612 N36612 0 diode
R36613 N36612 N36613 10
D36613 N36613 0 diode
R36614 N36613 N36614 10
D36614 N36614 0 diode
R36615 N36614 N36615 10
D36615 N36615 0 diode
R36616 N36615 N36616 10
D36616 N36616 0 diode
R36617 N36616 N36617 10
D36617 N36617 0 diode
R36618 N36617 N36618 10
D36618 N36618 0 diode
R36619 N36618 N36619 10
D36619 N36619 0 diode
R36620 N36619 N36620 10
D36620 N36620 0 diode
R36621 N36620 N36621 10
D36621 N36621 0 diode
R36622 N36621 N36622 10
D36622 N36622 0 diode
R36623 N36622 N36623 10
D36623 N36623 0 diode
R36624 N36623 N36624 10
D36624 N36624 0 diode
R36625 N36624 N36625 10
D36625 N36625 0 diode
R36626 N36625 N36626 10
D36626 N36626 0 diode
R36627 N36626 N36627 10
D36627 N36627 0 diode
R36628 N36627 N36628 10
D36628 N36628 0 diode
R36629 N36628 N36629 10
D36629 N36629 0 diode
R36630 N36629 N36630 10
D36630 N36630 0 diode
R36631 N36630 N36631 10
D36631 N36631 0 diode
R36632 N36631 N36632 10
D36632 N36632 0 diode
R36633 N36632 N36633 10
D36633 N36633 0 diode
R36634 N36633 N36634 10
D36634 N36634 0 diode
R36635 N36634 N36635 10
D36635 N36635 0 diode
R36636 N36635 N36636 10
D36636 N36636 0 diode
R36637 N36636 N36637 10
D36637 N36637 0 diode
R36638 N36637 N36638 10
D36638 N36638 0 diode
R36639 N36638 N36639 10
D36639 N36639 0 diode
R36640 N36639 N36640 10
D36640 N36640 0 diode
R36641 N36640 N36641 10
D36641 N36641 0 diode
R36642 N36641 N36642 10
D36642 N36642 0 diode
R36643 N36642 N36643 10
D36643 N36643 0 diode
R36644 N36643 N36644 10
D36644 N36644 0 diode
R36645 N36644 N36645 10
D36645 N36645 0 diode
R36646 N36645 N36646 10
D36646 N36646 0 diode
R36647 N36646 N36647 10
D36647 N36647 0 diode
R36648 N36647 N36648 10
D36648 N36648 0 diode
R36649 N36648 N36649 10
D36649 N36649 0 diode
R36650 N36649 N36650 10
D36650 N36650 0 diode
R36651 N36650 N36651 10
D36651 N36651 0 diode
R36652 N36651 N36652 10
D36652 N36652 0 diode
R36653 N36652 N36653 10
D36653 N36653 0 diode
R36654 N36653 N36654 10
D36654 N36654 0 diode
R36655 N36654 N36655 10
D36655 N36655 0 diode
R36656 N36655 N36656 10
D36656 N36656 0 diode
R36657 N36656 N36657 10
D36657 N36657 0 diode
R36658 N36657 N36658 10
D36658 N36658 0 diode
R36659 N36658 N36659 10
D36659 N36659 0 diode
R36660 N36659 N36660 10
D36660 N36660 0 diode
R36661 N36660 N36661 10
D36661 N36661 0 diode
R36662 N36661 N36662 10
D36662 N36662 0 diode
R36663 N36662 N36663 10
D36663 N36663 0 diode
R36664 N36663 N36664 10
D36664 N36664 0 diode
R36665 N36664 N36665 10
D36665 N36665 0 diode
R36666 N36665 N36666 10
D36666 N36666 0 diode
R36667 N36666 N36667 10
D36667 N36667 0 diode
R36668 N36667 N36668 10
D36668 N36668 0 diode
R36669 N36668 N36669 10
D36669 N36669 0 diode
R36670 N36669 N36670 10
D36670 N36670 0 diode
R36671 N36670 N36671 10
D36671 N36671 0 diode
R36672 N36671 N36672 10
D36672 N36672 0 diode
R36673 N36672 N36673 10
D36673 N36673 0 diode
R36674 N36673 N36674 10
D36674 N36674 0 diode
R36675 N36674 N36675 10
D36675 N36675 0 diode
R36676 N36675 N36676 10
D36676 N36676 0 diode
R36677 N36676 N36677 10
D36677 N36677 0 diode
R36678 N36677 N36678 10
D36678 N36678 0 diode
R36679 N36678 N36679 10
D36679 N36679 0 diode
R36680 N36679 N36680 10
D36680 N36680 0 diode
R36681 N36680 N36681 10
D36681 N36681 0 diode
R36682 N36681 N36682 10
D36682 N36682 0 diode
R36683 N36682 N36683 10
D36683 N36683 0 diode
R36684 N36683 N36684 10
D36684 N36684 0 diode
R36685 N36684 N36685 10
D36685 N36685 0 diode
R36686 N36685 N36686 10
D36686 N36686 0 diode
R36687 N36686 N36687 10
D36687 N36687 0 diode
R36688 N36687 N36688 10
D36688 N36688 0 diode
R36689 N36688 N36689 10
D36689 N36689 0 diode
R36690 N36689 N36690 10
D36690 N36690 0 diode
R36691 N36690 N36691 10
D36691 N36691 0 diode
R36692 N36691 N36692 10
D36692 N36692 0 diode
R36693 N36692 N36693 10
D36693 N36693 0 diode
R36694 N36693 N36694 10
D36694 N36694 0 diode
R36695 N36694 N36695 10
D36695 N36695 0 diode
R36696 N36695 N36696 10
D36696 N36696 0 diode
R36697 N36696 N36697 10
D36697 N36697 0 diode
R36698 N36697 N36698 10
D36698 N36698 0 diode
R36699 N36698 N36699 10
D36699 N36699 0 diode
R36700 N36699 N36700 10
D36700 N36700 0 diode
R36701 N36700 N36701 10
D36701 N36701 0 diode
R36702 N36701 N36702 10
D36702 N36702 0 diode
R36703 N36702 N36703 10
D36703 N36703 0 diode
R36704 N36703 N36704 10
D36704 N36704 0 diode
R36705 N36704 N36705 10
D36705 N36705 0 diode
R36706 N36705 N36706 10
D36706 N36706 0 diode
R36707 N36706 N36707 10
D36707 N36707 0 diode
R36708 N36707 N36708 10
D36708 N36708 0 diode
R36709 N36708 N36709 10
D36709 N36709 0 diode
R36710 N36709 N36710 10
D36710 N36710 0 diode
R36711 N36710 N36711 10
D36711 N36711 0 diode
R36712 N36711 N36712 10
D36712 N36712 0 diode
R36713 N36712 N36713 10
D36713 N36713 0 diode
R36714 N36713 N36714 10
D36714 N36714 0 diode
R36715 N36714 N36715 10
D36715 N36715 0 diode
R36716 N36715 N36716 10
D36716 N36716 0 diode
R36717 N36716 N36717 10
D36717 N36717 0 diode
R36718 N36717 N36718 10
D36718 N36718 0 diode
R36719 N36718 N36719 10
D36719 N36719 0 diode
R36720 N36719 N36720 10
D36720 N36720 0 diode
R36721 N36720 N36721 10
D36721 N36721 0 diode
R36722 N36721 N36722 10
D36722 N36722 0 diode
R36723 N36722 N36723 10
D36723 N36723 0 diode
R36724 N36723 N36724 10
D36724 N36724 0 diode
R36725 N36724 N36725 10
D36725 N36725 0 diode
R36726 N36725 N36726 10
D36726 N36726 0 diode
R36727 N36726 N36727 10
D36727 N36727 0 diode
R36728 N36727 N36728 10
D36728 N36728 0 diode
R36729 N36728 N36729 10
D36729 N36729 0 diode
R36730 N36729 N36730 10
D36730 N36730 0 diode
R36731 N36730 N36731 10
D36731 N36731 0 diode
R36732 N36731 N36732 10
D36732 N36732 0 diode
R36733 N36732 N36733 10
D36733 N36733 0 diode
R36734 N36733 N36734 10
D36734 N36734 0 diode
R36735 N36734 N36735 10
D36735 N36735 0 diode
R36736 N36735 N36736 10
D36736 N36736 0 diode
R36737 N36736 N36737 10
D36737 N36737 0 diode
R36738 N36737 N36738 10
D36738 N36738 0 diode
R36739 N36738 N36739 10
D36739 N36739 0 diode
R36740 N36739 N36740 10
D36740 N36740 0 diode
R36741 N36740 N36741 10
D36741 N36741 0 diode
R36742 N36741 N36742 10
D36742 N36742 0 diode
R36743 N36742 N36743 10
D36743 N36743 0 diode
R36744 N36743 N36744 10
D36744 N36744 0 diode
R36745 N36744 N36745 10
D36745 N36745 0 diode
R36746 N36745 N36746 10
D36746 N36746 0 diode
R36747 N36746 N36747 10
D36747 N36747 0 diode
R36748 N36747 N36748 10
D36748 N36748 0 diode
R36749 N36748 N36749 10
D36749 N36749 0 diode
R36750 N36749 N36750 10
D36750 N36750 0 diode
R36751 N36750 N36751 10
D36751 N36751 0 diode
R36752 N36751 N36752 10
D36752 N36752 0 diode
R36753 N36752 N36753 10
D36753 N36753 0 diode
R36754 N36753 N36754 10
D36754 N36754 0 diode
R36755 N36754 N36755 10
D36755 N36755 0 diode
R36756 N36755 N36756 10
D36756 N36756 0 diode
R36757 N36756 N36757 10
D36757 N36757 0 diode
R36758 N36757 N36758 10
D36758 N36758 0 diode
R36759 N36758 N36759 10
D36759 N36759 0 diode
R36760 N36759 N36760 10
D36760 N36760 0 diode
R36761 N36760 N36761 10
D36761 N36761 0 diode
R36762 N36761 N36762 10
D36762 N36762 0 diode
R36763 N36762 N36763 10
D36763 N36763 0 diode
R36764 N36763 N36764 10
D36764 N36764 0 diode
R36765 N36764 N36765 10
D36765 N36765 0 diode
R36766 N36765 N36766 10
D36766 N36766 0 diode
R36767 N36766 N36767 10
D36767 N36767 0 diode
R36768 N36767 N36768 10
D36768 N36768 0 diode
R36769 N36768 N36769 10
D36769 N36769 0 diode
R36770 N36769 N36770 10
D36770 N36770 0 diode
R36771 N36770 N36771 10
D36771 N36771 0 diode
R36772 N36771 N36772 10
D36772 N36772 0 diode
R36773 N36772 N36773 10
D36773 N36773 0 diode
R36774 N36773 N36774 10
D36774 N36774 0 diode
R36775 N36774 N36775 10
D36775 N36775 0 diode
R36776 N36775 N36776 10
D36776 N36776 0 diode
R36777 N36776 N36777 10
D36777 N36777 0 diode
R36778 N36777 N36778 10
D36778 N36778 0 diode
R36779 N36778 N36779 10
D36779 N36779 0 diode
R36780 N36779 N36780 10
D36780 N36780 0 diode
R36781 N36780 N36781 10
D36781 N36781 0 diode
R36782 N36781 N36782 10
D36782 N36782 0 diode
R36783 N36782 N36783 10
D36783 N36783 0 diode
R36784 N36783 N36784 10
D36784 N36784 0 diode
R36785 N36784 N36785 10
D36785 N36785 0 diode
R36786 N36785 N36786 10
D36786 N36786 0 diode
R36787 N36786 N36787 10
D36787 N36787 0 diode
R36788 N36787 N36788 10
D36788 N36788 0 diode
R36789 N36788 N36789 10
D36789 N36789 0 diode
R36790 N36789 N36790 10
D36790 N36790 0 diode
R36791 N36790 N36791 10
D36791 N36791 0 diode
R36792 N36791 N36792 10
D36792 N36792 0 diode
R36793 N36792 N36793 10
D36793 N36793 0 diode
R36794 N36793 N36794 10
D36794 N36794 0 diode
R36795 N36794 N36795 10
D36795 N36795 0 diode
R36796 N36795 N36796 10
D36796 N36796 0 diode
R36797 N36796 N36797 10
D36797 N36797 0 diode
R36798 N36797 N36798 10
D36798 N36798 0 diode
R36799 N36798 N36799 10
D36799 N36799 0 diode
R36800 N36799 N36800 10
D36800 N36800 0 diode
R36801 N36800 N36801 10
D36801 N36801 0 diode
R36802 N36801 N36802 10
D36802 N36802 0 diode
R36803 N36802 N36803 10
D36803 N36803 0 diode
R36804 N36803 N36804 10
D36804 N36804 0 diode
R36805 N36804 N36805 10
D36805 N36805 0 diode
R36806 N36805 N36806 10
D36806 N36806 0 diode
R36807 N36806 N36807 10
D36807 N36807 0 diode
R36808 N36807 N36808 10
D36808 N36808 0 diode
R36809 N36808 N36809 10
D36809 N36809 0 diode
R36810 N36809 N36810 10
D36810 N36810 0 diode
R36811 N36810 N36811 10
D36811 N36811 0 diode
R36812 N36811 N36812 10
D36812 N36812 0 diode
R36813 N36812 N36813 10
D36813 N36813 0 diode
R36814 N36813 N36814 10
D36814 N36814 0 diode
R36815 N36814 N36815 10
D36815 N36815 0 diode
R36816 N36815 N36816 10
D36816 N36816 0 diode
R36817 N36816 N36817 10
D36817 N36817 0 diode
R36818 N36817 N36818 10
D36818 N36818 0 diode
R36819 N36818 N36819 10
D36819 N36819 0 diode
R36820 N36819 N36820 10
D36820 N36820 0 diode
R36821 N36820 N36821 10
D36821 N36821 0 diode
R36822 N36821 N36822 10
D36822 N36822 0 diode
R36823 N36822 N36823 10
D36823 N36823 0 diode
R36824 N36823 N36824 10
D36824 N36824 0 diode
R36825 N36824 N36825 10
D36825 N36825 0 diode
R36826 N36825 N36826 10
D36826 N36826 0 diode
R36827 N36826 N36827 10
D36827 N36827 0 diode
R36828 N36827 N36828 10
D36828 N36828 0 diode
R36829 N36828 N36829 10
D36829 N36829 0 diode
R36830 N36829 N36830 10
D36830 N36830 0 diode
R36831 N36830 N36831 10
D36831 N36831 0 diode
R36832 N36831 N36832 10
D36832 N36832 0 diode
R36833 N36832 N36833 10
D36833 N36833 0 diode
R36834 N36833 N36834 10
D36834 N36834 0 diode
R36835 N36834 N36835 10
D36835 N36835 0 diode
R36836 N36835 N36836 10
D36836 N36836 0 diode
R36837 N36836 N36837 10
D36837 N36837 0 diode
R36838 N36837 N36838 10
D36838 N36838 0 diode
R36839 N36838 N36839 10
D36839 N36839 0 diode
R36840 N36839 N36840 10
D36840 N36840 0 diode
R36841 N36840 N36841 10
D36841 N36841 0 diode
R36842 N36841 N36842 10
D36842 N36842 0 diode
R36843 N36842 N36843 10
D36843 N36843 0 diode
R36844 N36843 N36844 10
D36844 N36844 0 diode
R36845 N36844 N36845 10
D36845 N36845 0 diode
R36846 N36845 N36846 10
D36846 N36846 0 diode
R36847 N36846 N36847 10
D36847 N36847 0 diode
R36848 N36847 N36848 10
D36848 N36848 0 diode
R36849 N36848 N36849 10
D36849 N36849 0 diode
R36850 N36849 N36850 10
D36850 N36850 0 diode
R36851 N36850 N36851 10
D36851 N36851 0 diode
R36852 N36851 N36852 10
D36852 N36852 0 diode
R36853 N36852 N36853 10
D36853 N36853 0 diode
R36854 N36853 N36854 10
D36854 N36854 0 diode
R36855 N36854 N36855 10
D36855 N36855 0 diode
R36856 N36855 N36856 10
D36856 N36856 0 diode
R36857 N36856 N36857 10
D36857 N36857 0 diode
R36858 N36857 N36858 10
D36858 N36858 0 diode
R36859 N36858 N36859 10
D36859 N36859 0 diode
R36860 N36859 N36860 10
D36860 N36860 0 diode
R36861 N36860 N36861 10
D36861 N36861 0 diode
R36862 N36861 N36862 10
D36862 N36862 0 diode
R36863 N36862 N36863 10
D36863 N36863 0 diode
R36864 N36863 N36864 10
D36864 N36864 0 diode
R36865 N36864 N36865 10
D36865 N36865 0 diode
R36866 N36865 N36866 10
D36866 N36866 0 diode
R36867 N36866 N36867 10
D36867 N36867 0 diode
R36868 N36867 N36868 10
D36868 N36868 0 diode
R36869 N36868 N36869 10
D36869 N36869 0 diode
R36870 N36869 N36870 10
D36870 N36870 0 diode
R36871 N36870 N36871 10
D36871 N36871 0 diode
R36872 N36871 N36872 10
D36872 N36872 0 diode
R36873 N36872 N36873 10
D36873 N36873 0 diode
R36874 N36873 N36874 10
D36874 N36874 0 diode
R36875 N36874 N36875 10
D36875 N36875 0 diode
R36876 N36875 N36876 10
D36876 N36876 0 diode
R36877 N36876 N36877 10
D36877 N36877 0 diode
R36878 N36877 N36878 10
D36878 N36878 0 diode
R36879 N36878 N36879 10
D36879 N36879 0 diode
R36880 N36879 N36880 10
D36880 N36880 0 diode
R36881 N36880 N36881 10
D36881 N36881 0 diode
R36882 N36881 N36882 10
D36882 N36882 0 diode
R36883 N36882 N36883 10
D36883 N36883 0 diode
R36884 N36883 N36884 10
D36884 N36884 0 diode
R36885 N36884 N36885 10
D36885 N36885 0 diode
R36886 N36885 N36886 10
D36886 N36886 0 diode
R36887 N36886 N36887 10
D36887 N36887 0 diode
R36888 N36887 N36888 10
D36888 N36888 0 diode
R36889 N36888 N36889 10
D36889 N36889 0 diode
R36890 N36889 N36890 10
D36890 N36890 0 diode
R36891 N36890 N36891 10
D36891 N36891 0 diode
R36892 N36891 N36892 10
D36892 N36892 0 diode
R36893 N36892 N36893 10
D36893 N36893 0 diode
R36894 N36893 N36894 10
D36894 N36894 0 diode
R36895 N36894 N36895 10
D36895 N36895 0 diode
R36896 N36895 N36896 10
D36896 N36896 0 diode
R36897 N36896 N36897 10
D36897 N36897 0 diode
R36898 N36897 N36898 10
D36898 N36898 0 diode
R36899 N36898 N36899 10
D36899 N36899 0 diode
R36900 N36899 N36900 10
D36900 N36900 0 diode
R36901 N36900 N36901 10
D36901 N36901 0 diode
R36902 N36901 N36902 10
D36902 N36902 0 diode
R36903 N36902 N36903 10
D36903 N36903 0 diode
R36904 N36903 N36904 10
D36904 N36904 0 diode
R36905 N36904 N36905 10
D36905 N36905 0 diode
R36906 N36905 N36906 10
D36906 N36906 0 diode
R36907 N36906 N36907 10
D36907 N36907 0 diode
R36908 N36907 N36908 10
D36908 N36908 0 diode
R36909 N36908 N36909 10
D36909 N36909 0 diode
R36910 N36909 N36910 10
D36910 N36910 0 diode
R36911 N36910 N36911 10
D36911 N36911 0 diode
R36912 N36911 N36912 10
D36912 N36912 0 diode
R36913 N36912 N36913 10
D36913 N36913 0 diode
R36914 N36913 N36914 10
D36914 N36914 0 diode
R36915 N36914 N36915 10
D36915 N36915 0 diode
R36916 N36915 N36916 10
D36916 N36916 0 diode
R36917 N36916 N36917 10
D36917 N36917 0 diode
R36918 N36917 N36918 10
D36918 N36918 0 diode
R36919 N36918 N36919 10
D36919 N36919 0 diode
R36920 N36919 N36920 10
D36920 N36920 0 diode
R36921 N36920 N36921 10
D36921 N36921 0 diode
R36922 N36921 N36922 10
D36922 N36922 0 diode
R36923 N36922 N36923 10
D36923 N36923 0 diode
R36924 N36923 N36924 10
D36924 N36924 0 diode
R36925 N36924 N36925 10
D36925 N36925 0 diode
R36926 N36925 N36926 10
D36926 N36926 0 diode
R36927 N36926 N36927 10
D36927 N36927 0 diode
R36928 N36927 N36928 10
D36928 N36928 0 diode
R36929 N36928 N36929 10
D36929 N36929 0 diode
R36930 N36929 N36930 10
D36930 N36930 0 diode
R36931 N36930 N36931 10
D36931 N36931 0 diode
R36932 N36931 N36932 10
D36932 N36932 0 diode
R36933 N36932 N36933 10
D36933 N36933 0 diode
R36934 N36933 N36934 10
D36934 N36934 0 diode
R36935 N36934 N36935 10
D36935 N36935 0 diode
R36936 N36935 N36936 10
D36936 N36936 0 diode
R36937 N36936 N36937 10
D36937 N36937 0 diode
R36938 N36937 N36938 10
D36938 N36938 0 diode
R36939 N36938 N36939 10
D36939 N36939 0 diode
R36940 N36939 N36940 10
D36940 N36940 0 diode
R36941 N36940 N36941 10
D36941 N36941 0 diode
R36942 N36941 N36942 10
D36942 N36942 0 diode
R36943 N36942 N36943 10
D36943 N36943 0 diode
R36944 N36943 N36944 10
D36944 N36944 0 diode
R36945 N36944 N36945 10
D36945 N36945 0 diode
R36946 N36945 N36946 10
D36946 N36946 0 diode
R36947 N36946 N36947 10
D36947 N36947 0 diode
R36948 N36947 N36948 10
D36948 N36948 0 diode
R36949 N36948 N36949 10
D36949 N36949 0 diode
R36950 N36949 N36950 10
D36950 N36950 0 diode
R36951 N36950 N36951 10
D36951 N36951 0 diode
R36952 N36951 N36952 10
D36952 N36952 0 diode
R36953 N36952 N36953 10
D36953 N36953 0 diode
R36954 N36953 N36954 10
D36954 N36954 0 diode
R36955 N36954 N36955 10
D36955 N36955 0 diode
R36956 N36955 N36956 10
D36956 N36956 0 diode
R36957 N36956 N36957 10
D36957 N36957 0 diode
R36958 N36957 N36958 10
D36958 N36958 0 diode
R36959 N36958 N36959 10
D36959 N36959 0 diode
R36960 N36959 N36960 10
D36960 N36960 0 diode
R36961 N36960 N36961 10
D36961 N36961 0 diode
R36962 N36961 N36962 10
D36962 N36962 0 diode
R36963 N36962 N36963 10
D36963 N36963 0 diode
R36964 N36963 N36964 10
D36964 N36964 0 diode
R36965 N36964 N36965 10
D36965 N36965 0 diode
R36966 N36965 N36966 10
D36966 N36966 0 diode
R36967 N36966 N36967 10
D36967 N36967 0 diode
R36968 N36967 N36968 10
D36968 N36968 0 diode
R36969 N36968 N36969 10
D36969 N36969 0 diode
R36970 N36969 N36970 10
D36970 N36970 0 diode
R36971 N36970 N36971 10
D36971 N36971 0 diode
R36972 N36971 N36972 10
D36972 N36972 0 diode
R36973 N36972 N36973 10
D36973 N36973 0 diode
R36974 N36973 N36974 10
D36974 N36974 0 diode
R36975 N36974 N36975 10
D36975 N36975 0 diode
R36976 N36975 N36976 10
D36976 N36976 0 diode
R36977 N36976 N36977 10
D36977 N36977 0 diode
R36978 N36977 N36978 10
D36978 N36978 0 diode
R36979 N36978 N36979 10
D36979 N36979 0 diode
R36980 N36979 N36980 10
D36980 N36980 0 diode
R36981 N36980 N36981 10
D36981 N36981 0 diode
R36982 N36981 N36982 10
D36982 N36982 0 diode
R36983 N36982 N36983 10
D36983 N36983 0 diode
R36984 N36983 N36984 10
D36984 N36984 0 diode
R36985 N36984 N36985 10
D36985 N36985 0 diode
R36986 N36985 N36986 10
D36986 N36986 0 diode
R36987 N36986 N36987 10
D36987 N36987 0 diode
R36988 N36987 N36988 10
D36988 N36988 0 diode
R36989 N36988 N36989 10
D36989 N36989 0 diode
R36990 N36989 N36990 10
D36990 N36990 0 diode
R36991 N36990 N36991 10
D36991 N36991 0 diode
R36992 N36991 N36992 10
D36992 N36992 0 diode
R36993 N36992 N36993 10
D36993 N36993 0 diode
R36994 N36993 N36994 10
D36994 N36994 0 diode
R36995 N36994 N36995 10
D36995 N36995 0 diode
R36996 N36995 N36996 10
D36996 N36996 0 diode
R36997 N36996 N36997 10
D36997 N36997 0 diode
R36998 N36997 N36998 10
D36998 N36998 0 diode
R36999 N36998 N36999 10
D36999 N36999 0 diode
R37000 N36999 N37000 10
D37000 N37000 0 diode
R37001 N37000 N37001 10
D37001 N37001 0 diode
R37002 N37001 N37002 10
D37002 N37002 0 diode
R37003 N37002 N37003 10
D37003 N37003 0 diode
R37004 N37003 N37004 10
D37004 N37004 0 diode
R37005 N37004 N37005 10
D37005 N37005 0 diode
R37006 N37005 N37006 10
D37006 N37006 0 diode
R37007 N37006 N37007 10
D37007 N37007 0 diode
R37008 N37007 N37008 10
D37008 N37008 0 diode
R37009 N37008 N37009 10
D37009 N37009 0 diode
R37010 N37009 N37010 10
D37010 N37010 0 diode
R37011 N37010 N37011 10
D37011 N37011 0 diode
R37012 N37011 N37012 10
D37012 N37012 0 diode
R37013 N37012 N37013 10
D37013 N37013 0 diode
R37014 N37013 N37014 10
D37014 N37014 0 diode
R37015 N37014 N37015 10
D37015 N37015 0 diode
R37016 N37015 N37016 10
D37016 N37016 0 diode
R37017 N37016 N37017 10
D37017 N37017 0 diode
R37018 N37017 N37018 10
D37018 N37018 0 diode
R37019 N37018 N37019 10
D37019 N37019 0 diode
R37020 N37019 N37020 10
D37020 N37020 0 diode
R37021 N37020 N37021 10
D37021 N37021 0 diode
R37022 N37021 N37022 10
D37022 N37022 0 diode
R37023 N37022 N37023 10
D37023 N37023 0 diode
R37024 N37023 N37024 10
D37024 N37024 0 diode
R37025 N37024 N37025 10
D37025 N37025 0 diode
R37026 N37025 N37026 10
D37026 N37026 0 diode
R37027 N37026 N37027 10
D37027 N37027 0 diode
R37028 N37027 N37028 10
D37028 N37028 0 diode
R37029 N37028 N37029 10
D37029 N37029 0 diode
R37030 N37029 N37030 10
D37030 N37030 0 diode
R37031 N37030 N37031 10
D37031 N37031 0 diode
R37032 N37031 N37032 10
D37032 N37032 0 diode
R37033 N37032 N37033 10
D37033 N37033 0 diode
R37034 N37033 N37034 10
D37034 N37034 0 diode
R37035 N37034 N37035 10
D37035 N37035 0 diode
R37036 N37035 N37036 10
D37036 N37036 0 diode
R37037 N37036 N37037 10
D37037 N37037 0 diode
R37038 N37037 N37038 10
D37038 N37038 0 diode
R37039 N37038 N37039 10
D37039 N37039 0 diode
R37040 N37039 N37040 10
D37040 N37040 0 diode
R37041 N37040 N37041 10
D37041 N37041 0 diode
R37042 N37041 N37042 10
D37042 N37042 0 diode
R37043 N37042 N37043 10
D37043 N37043 0 diode
R37044 N37043 N37044 10
D37044 N37044 0 diode
R37045 N37044 N37045 10
D37045 N37045 0 diode
R37046 N37045 N37046 10
D37046 N37046 0 diode
R37047 N37046 N37047 10
D37047 N37047 0 diode
R37048 N37047 N37048 10
D37048 N37048 0 diode
R37049 N37048 N37049 10
D37049 N37049 0 diode
R37050 N37049 N37050 10
D37050 N37050 0 diode
R37051 N37050 N37051 10
D37051 N37051 0 diode
R37052 N37051 N37052 10
D37052 N37052 0 diode
R37053 N37052 N37053 10
D37053 N37053 0 diode
R37054 N37053 N37054 10
D37054 N37054 0 diode
R37055 N37054 N37055 10
D37055 N37055 0 diode
R37056 N37055 N37056 10
D37056 N37056 0 diode
R37057 N37056 N37057 10
D37057 N37057 0 diode
R37058 N37057 N37058 10
D37058 N37058 0 diode
R37059 N37058 N37059 10
D37059 N37059 0 diode
R37060 N37059 N37060 10
D37060 N37060 0 diode
R37061 N37060 N37061 10
D37061 N37061 0 diode
R37062 N37061 N37062 10
D37062 N37062 0 diode
R37063 N37062 N37063 10
D37063 N37063 0 diode
R37064 N37063 N37064 10
D37064 N37064 0 diode
R37065 N37064 N37065 10
D37065 N37065 0 diode
R37066 N37065 N37066 10
D37066 N37066 0 diode
R37067 N37066 N37067 10
D37067 N37067 0 diode
R37068 N37067 N37068 10
D37068 N37068 0 diode
R37069 N37068 N37069 10
D37069 N37069 0 diode
R37070 N37069 N37070 10
D37070 N37070 0 diode
R37071 N37070 N37071 10
D37071 N37071 0 diode
R37072 N37071 N37072 10
D37072 N37072 0 diode
R37073 N37072 N37073 10
D37073 N37073 0 diode
R37074 N37073 N37074 10
D37074 N37074 0 diode
R37075 N37074 N37075 10
D37075 N37075 0 diode
R37076 N37075 N37076 10
D37076 N37076 0 diode
R37077 N37076 N37077 10
D37077 N37077 0 diode
R37078 N37077 N37078 10
D37078 N37078 0 diode
R37079 N37078 N37079 10
D37079 N37079 0 diode
R37080 N37079 N37080 10
D37080 N37080 0 diode
R37081 N37080 N37081 10
D37081 N37081 0 diode
R37082 N37081 N37082 10
D37082 N37082 0 diode
R37083 N37082 N37083 10
D37083 N37083 0 diode
R37084 N37083 N37084 10
D37084 N37084 0 diode
R37085 N37084 N37085 10
D37085 N37085 0 diode
R37086 N37085 N37086 10
D37086 N37086 0 diode
R37087 N37086 N37087 10
D37087 N37087 0 diode
R37088 N37087 N37088 10
D37088 N37088 0 diode
R37089 N37088 N37089 10
D37089 N37089 0 diode
R37090 N37089 N37090 10
D37090 N37090 0 diode
R37091 N37090 N37091 10
D37091 N37091 0 diode
R37092 N37091 N37092 10
D37092 N37092 0 diode
R37093 N37092 N37093 10
D37093 N37093 0 diode
R37094 N37093 N37094 10
D37094 N37094 0 diode
R37095 N37094 N37095 10
D37095 N37095 0 diode
R37096 N37095 N37096 10
D37096 N37096 0 diode
R37097 N37096 N37097 10
D37097 N37097 0 diode
R37098 N37097 N37098 10
D37098 N37098 0 diode
R37099 N37098 N37099 10
D37099 N37099 0 diode
R37100 N37099 N37100 10
D37100 N37100 0 diode
R37101 N37100 N37101 10
D37101 N37101 0 diode
R37102 N37101 N37102 10
D37102 N37102 0 diode
R37103 N37102 N37103 10
D37103 N37103 0 diode
R37104 N37103 N37104 10
D37104 N37104 0 diode
R37105 N37104 N37105 10
D37105 N37105 0 diode
R37106 N37105 N37106 10
D37106 N37106 0 diode
R37107 N37106 N37107 10
D37107 N37107 0 diode
R37108 N37107 N37108 10
D37108 N37108 0 diode
R37109 N37108 N37109 10
D37109 N37109 0 diode
R37110 N37109 N37110 10
D37110 N37110 0 diode
R37111 N37110 N37111 10
D37111 N37111 0 diode
R37112 N37111 N37112 10
D37112 N37112 0 diode
R37113 N37112 N37113 10
D37113 N37113 0 diode
R37114 N37113 N37114 10
D37114 N37114 0 diode
R37115 N37114 N37115 10
D37115 N37115 0 diode
R37116 N37115 N37116 10
D37116 N37116 0 diode
R37117 N37116 N37117 10
D37117 N37117 0 diode
R37118 N37117 N37118 10
D37118 N37118 0 diode
R37119 N37118 N37119 10
D37119 N37119 0 diode
R37120 N37119 N37120 10
D37120 N37120 0 diode
R37121 N37120 N37121 10
D37121 N37121 0 diode
R37122 N37121 N37122 10
D37122 N37122 0 diode
R37123 N37122 N37123 10
D37123 N37123 0 diode
R37124 N37123 N37124 10
D37124 N37124 0 diode
R37125 N37124 N37125 10
D37125 N37125 0 diode
R37126 N37125 N37126 10
D37126 N37126 0 diode
R37127 N37126 N37127 10
D37127 N37127 0 diode
R37128 N37127 N37128 10
D37128 N37128 0 diode
R37129 N37128 N37129 10
D37129 N37129 0 diode
R37130 N37129 N37130 10
D37130 N37130 0 diode
R37131 N37130 N37131 10
D37131 N37131 0 diode
R37132 N37131 N37132 10
D37132 N37132 0 diode
R37133 N37132 N37133 10
D37133 N37133 0 diode
R37134 N37133 N37134 10
D37134 N37134 0 diode
R37135 N37134 N37135 10
D37135 N37135 0 diode
R37136 N37135 N37136 10
D37136 N37136 0 diode
R37137 N37136 N37137 10
D37137 N37137 0 diode
R37138 N37137 N37138 10
D37138 N37138 0 diode
R37139 N37138 N37139 10
D37139 N37139 0 diode
R37140 N37139 N37140 10
D37140 N37140 0 diode
R37141 N37140 N37141 10
D37141 N37141 0 diode
R37142 N37141 N37142 10
D37142 N37142 0 diode
R37143 N37142 N37143 10
D37143 N37143 0 diode
R37144 N37143 N37144 10
D37144 N37144 0 diode
R37145 N37144 N37145 10
D37145 N37145 0 diode
R37146 N37145 N37146 10
D37146 N37146 0 diode
R37147 N37146 N37147 10
D37147 N37147 0 diode
R37148 N37147 N37148 10
D37148 N37148 0 diode
R37149 N37148 N37149 10
D37149 N37149 0 diode
R37150 N37149 N37150 10
D37150 N37150 0 diode
R37151 N37150 N37151 10
D37151 N37151 0 diode
R37152 N37151 N37152 10
D37152 N37152 0 diode
R37153 N37152 N37153 10
D37153 N37153 0 diode
R37154 N37153 N37154 10
D37154 N37154 0 diode
R37155 N37154 N37155 10
D37155 N37155 0 diode
R37156 N37155 N37156 10
D37156 N37156 0 diode
R37157 N37156 N37157 10
D37157 N37157 0 diode
R37158 N37157 N37158 10
D37158 N37158 0 diode
R37159 N37158 N37159 10
D37159 N37159 0 diode
R37160 N37159 N37160 10
D37160 N37160 0 diode
R37161 N37160 N37161 10
D37161 N37161 0 diode
R37162 N37161 N37162 10
D37162 N37162 0 diode
R37163 N37162 N37163 10
D37163 N37163 0 diode
R37164 N37163 N37164 10
D37164 N37164 0 diode
R37165 N37164 N37165 10
D37165 N37165 0 diode
R37166 N37165 N37166 10
D37166 N37166 0 diode
R37167 N37166 N37167 10
D37167 N37167 0 diode
R37168 N37167 N37168 10
D37168 N37168 0 diode
R37169 N37168 N37169 10
D37169 N37169 0 diode
R37170 N37169 N37170 10
D37170 N37170 0 diode
R37171 N37170 N37171 10
D37171 N37171 0 diode
R37172 N37171 N37172 10
D37172 N37172 0 diode
R37173 N37172 N37173 10
D37173 N37173 0 diode
R37174 N37173 N37174 10
D37174 N37174 0 diode
R37175 N37174 N37175 10
D37175 N37175 0 diode
R37176 N37175 N37176 10
D37176 N37176 0 diode
R37177 N37176 N37177 10
D37177 N37177 0 diode
R37178 N37177 N37178 10
D37178 N37178 0 diode
R37179 N37178 N37179 10
D37179 N37179 0 diode
R37180 N37179 N37180 10
D37180 N37180 0 diode
R37181 N37180 N37181 10
D37181 N37181 0 diode
R37182 N37181 N37182 10
D37182 N37182 0 diode
R37183 N37182 N37183 10
D37183 N37183 0 diode
R37184 N37183 N37184 10
D37184 N37184 0 diode
R37185 N37184 N37185 10
D37185 N37185 0 diode
R37186 N37185 N37186 10
D37186 N37186 0 diode
R37187 N37186 N37187 10
D37187 N37187 0 diode
R37188 N37187 N37188 10
D37188 N37188 0 diode
R37189 N37188 N37189 10
D37189 N37189 0 diode
R37190 N37189 N37190 10
D37190 N37190 0 diode
R37191 N37190 N37191 10
D37191 N37191 0 diode
R37192 N37191 N37192 10
D37192 N37192 0 diode
R37193 N37192 N37193 10
D37193 N37193 0 diode
R37194 N37193 N37194 10
D37194 N37194 0 diode
R37195 N37194 N37195 10
D37195 N37195 0 diode
R37196 N37195 N37196 10
D37196 N37196 0 diode
R37197 N37196 N37197 10
D37197 N37197 0 diode
R37198 N37197 N37198 10
D37198 N37198 0 diode
R37199 N37198 N37199 10
D37199 N37199 0 diode
R37200 N37199 N37200 10
D37200 N37200 0 diode
R37201 N37200 N37201 10
D37201 N37201 0 diode
R37202 N37201 N37202 10
D37202 N37202 0 diode
R37203 N37202 N37203 10
D37203 N37203 0 diode
R37204 N37203 N37204 10
D37204 N37204 0 diode
R37205 N37204 N37205 10
D37205 N37205 0 diode
R37206 N37205 N37206 10
D37206 N37206 0 diode
R37207 N37206 N37207 10
D37207 N37207 0 diode
R37208 N37207 N37208 10
D37208 N37208 0 diode
R37209 N37208 N37209 10
D37209 N37209 0 diode
R37210 N37209 N37210 10
D37210 N37210 0 diode
R37211 N37210 N37211 10
D37211 N37211 0 diode
R37212 N37211 N37212 10
D37212 N37212 0 diode
R37213 N37212 N37213 10
D37213 N37213 0 diode
R37214 N37213 N37214 10
D37214 N37214 0 diode
R37215 N37214 N37215 10
D37215 N37215 0 diode
R37216 N37215 N37216 10
D37216 N37216 0 diode
R37217 N37216 N37217 10
D37217 N37217 0 diode
R37218 N37217 N37218 10
D37218 N37218 0 diode
R37219 N37218 N37219 10
D37219 N37219 0 diode
R37220 N37219 N37220 10
D37220 N37220 0 diode
R37221 N37220 N37221 10
D37221 N37221 0 diode
R37222 N37221 N37222 10
D37222 N37222 0 diode
R37223 N37222 N37223 10
D37223 N37223 0 diode
R37224 N37223 N37224 10
D37224 N37224 0 diode
R37225 N37224 N37225 10
D37225 N37225 0 diode
R37226 N37225 N37226 10
D37226 N37226 0 diode
R37227 N37226 N37227 10
D37227 N37227 0 diode
R37228 N37227 N37228 10
D37228 N37228 0 diode
R37229 N37228 N37229 10
D37229 N37229 0 diode
R37230 N37229 N37230 10
D37230 N37230 0 diode
R37231 N37230 N37231 10
D37231 N37231 0 diode
R37232 N37231 N37232 10
D37232 N37232 0 diode
R37233 N37232 N37233 10
D37233 N37233 0 diode
R37234 N37233 N37234 10
D37234 N37234 0 diode
R37235 N37234 N37235 10
D37235 N37235 0 diode
R37236 N37235 N37236 10
D37236 N37236 0 diode
R37237 N37236 N37237 10
D37237 N37237 0 diode
R37238 N37237 N37238 10
D37238 N37238 0 diode
R37239 N37238 N37239 10
D37239 N37239 0 diode
R37240 N37239 N37240 10
D37240 N37240 0 diode
R37241 N37240 N37241 10
D37241 N37241 0 diode
R37242 N37241 N37242 10
D37242 N37242 0 diode
R37243 N37242 N37243 10
D37243 N37243 0 diode
R37244 N37243 N37244 10
D37244 N37244 0 diode
R37245 N37244 N37245 10
D37245 N37245 0 diode
R37246 N37245 N37246 10
D37246 N37246 0 diode
R37247 N37246 N37247 10
D37247 N37247 0 diode
R37248 N37247 N37248 10
D37248 N37248 0 diode
R37249 N37248 N37249 10
D37249 N37249 0 diode
R37250 N37249 N37250 10
D37250 N37250 0 diode
R37251 N37250 N37251 10
D37251 N37251 0 diode
R37252 N37251 N37252 10
D37252 N37252 0 diode
R37253 N37252 N37253 10
D37253 N37253 0 diode
R37254 N37253 N37254 10
D37254 N37254 0 diode
R37255 N37254 N37255 10
D37255 N37255 0 diode
R37256 N37255 N37256 10
D37256 N37256 0 diode
R37257 N37256 N37257 10
D37257 N37257 0 diode
R37258 N37257 N37258 10
D37258 N37258 0 diode
R37259 N37258 N37259 10
D37259 N37259 0 diode
R37260 N37259 N37260 10
D37260 N37260 0 diode
R37261 N37260 N37261 10
D37261 N37261 0 diode
R37262 N37261 N37262 10
D37262 N37262 0 diode
R37263 N37262 N37263 10
D37263 N37263 0 diode
R37264 N37263 N37264 10
D37264 N37264 0 diode
R37265 N37264 N37265 10
D37265 N37265 0 diode
R37266 N37265 N37266 10
D37266 N37266 0 diode
R37267 N37266 N37267 10
D37267 N37267 0 diode
R37268 N37267 N37268 10
D37268 N37268 0 diode
R37269 N37268 N37269 10
D37269 N37269 0 diode
R37270 N37269 N37270 10
D37270 N37270 0 diode
R37271 N37270 N37271 10
D37271 N37271 0 diode
R37272 N37271 N37272 10
D37272 N37272 0 diode
R37273 N37272 N37273 10
D37273 N37273 0 diode
R37274 N37273 N37274 10
D37274 N37274 0 diode
R37275 N37274 N37275 10
D37275 N37275 0 diode
R37276 N37275 N37276 10
D37276 N37276 0 diode
R37277 N37276 N37277 10
D37277 N37277 0 diode
R37278 N37277 N37278 10
D37278 N37278 0 diode
R37279 N37278 N37279 10
D37279 N37279 0 diode
R37280 N37279 N37280 10
D37280 N37280 0 diode
R37281 N37280 N37281 10
D37281 N37281 0 diode
R37282 N37281 N37282 10
D37282 N37282 0 diode
R37283 N37282 N37283 10
D37283 N37283 0 diode
R37284 N37283 N37284 10
D37284 N37284 0 diode
R37285 N37284 N37285 10
D37285 N37285 0 diode
R37286 N37285 N37286 10
D37286 N37286 0 diode
R37287 N37286 N37287 10
D37287 N37287 0 diode
R37288 N37287 N37288 10
D37288 N37288 0 diode
R37289 N37288 N37289 10
D37289 N37289 0 diode
R37290 N37289 N37290 10
D37290 N37290 0 diode
R37291 N37290 N37291 10
D37291 N37291 0 diode
R37292 N37291 N37292 10
D37292 N37292 0 diode
R37293 N37292 N37293 10
D37293 N37293 0 diode
R37294 N37293 N37294 10
D37294 N37294 0 diode
R37295 N37294 N37295 10
D37295 N37295 0 diode
R37296 N37295 N37296 10
D37296 N37296 0 diode
R37297 N37296 N37297 10
D37297 N37297 0 diode
R37298 N37297 N37298 10
D37298 N37298 0 diode
R37299 N37298 N37299 10
D37299 N37299 0 diode
R37300 N37299 N37300 10
D37300 N37300 0 diode
R37301 N37300 N37301 10
D37301 N37301 0 diode
R37302 N37301 N37302 10
D37302 N37302 0 diode
R37303 N37302 N37303 10
D37303 N37303 0 diode
R37304 N37303 N37304 10
D37304 N37304 0 diode
R37305 N37304 N37305 10
D37305 N37305 0 diode
R37306 N37305 N37306 10
D37306 N37306 0 diode
R37307 N37306 N37307 10
D37307 N37307 0 diode
R37308 N37307 N37308 10
D37308 N37308 0 diode
R37309 N37308 N37309 10
D37309 N37309 0 diode
R37310 N37309 N37310 10
D37310 N37310 0 diode
R37311 N37310 N37311 10
D37311 N37311 0 diode
R37312 N37311 N37312 10
D37312 N37312 0 diode
R37313 N37312 N37313 10
D37313 N37313 0 diode
R37314 N37313 N37314 10
D37314 N37314 0 diode
R37315 N37314 N37315 10
D37315 N37315 0 diode
R37316 N37315 N37316 10
D37316 N37316 0 diode
R37317 N37316 N37317 10
D37317 N37317 0 diode
R37318 N37317 N37318 10
D37318 N37318 0 diode
R37319 N37318 N37319 10
D37319 N37319 0 diode
R37320 N37319 N37320 10
D37320 N37320 0 diode
R37321 N37320 N37321 10
D37321 N37321 0 diode
R37322 N37321 N37322 10
D37322 N37322 0 diode
R37323 N37322 N37323 10
D37323 N37323 0 diode
R37324 N37323 N37324 10
D37324 N37324 0 diode
R37325 N37324 N37325 10
D37325 N37325 0 diode
R37326 N37325 N37326 10
D37326 N37326 0 diode
R37327 N37326 N37327 10
D37327 N37327 0 diode
R37328 N37327 N37328 10
D37328 N37328 0 diode
R37329 N37328 N37329 10
D37329 N37329 0 diode
R37330 N37329 N37330 10
D37330 N37330 0 diode
R37331 N37330 N37331 10
D37331 N37331 0 diode
R37332 N37331 N37332 10
D37332 N37332 0 diode
R37333 N37332 N37333 10
D37333 N37333 0 diode
R37334 N37333 N37334 10
D37334 N37334 0 diode
R37335 N37334 N37335 10
D37335 N37335 0 diode
R37336 N37335 N37336 10
D37336 N37336 0 diode
R37337 N37336 N37337 10
D37337 N37337 0 diode
R37338 N37337 N37338 10
D37338 N37338 0 diode
R37339 N37338 N37339 10
D37339 N37339 0 diode
R37340 N37339 N37340 10
D37340 N37340 0 diode
R37341 N37340 N37341 10
D37341 N37341 0 diode
R37342 N37341 N37342 10
D37342 N37342 0 diode
R37343 N37342 N37343 10
D37343 N37343 0 diode
R37344 N37343 N37344 10
D37344 N37344 0 diode
R37345 N37344 N37345 10
D37345 N37345 0 diode
R37346 N37345 N37346 10
D37346 N37346 0 diode
R37347 N37346 N37347 10
D37347 N37347 0 diode
R37348 N37347 N37348 10
D37348 N37348 0 diode
R37349 N37348 N37349 10
D37349 N37349 0 diode
R37350 N37349 N37350 10
D37350 N37350 0 diode
R37351 N37350 N37351 10
D37351 N37351 0 diode
R37352 N37351 N37352 10
D37352 N37352 0 diode
R37353 N37352 N37353 10
D37353 N37353 0 diode
R37354 N37353 N37354 10
D37354 N37354 0 diode
R37355 N37354 N37355 10
D37355 N37355 0 diode
R37356 N37355 N37356 10
D37356 N37356 0 diode
R37357 N37356 N37357 10
D37357 N37357 0 diode
R37358 N37357 N37358 10
D37358 N37358 0 diode
R37359 N37358 N37359 10
D37359 N37359 0 diode
R37360 N37359 N37360 10
D37360 N37360 0 diode
R37361 N37360 N37361 10
D37361 N37361 0 diode
R37362 N37361 N37362 10
D37362 N37362 0 diode
R37363 N37362 N37363 10
D37363 N37363 0 diode
R37364 N37363 N37364 10
D37364 N37364 0 diode
R37365 N37364 N37365 10
D37365 N37365 0 diode
R37366 N37365 N37366 10
D37366 N37366 0 diode
R37367 N37366 N37367 10
D37367 N37367 0 diode
R37368 N37367 N37368 10
D37368 N37368 0 diode
R37369 N37368 N37369 10
D37369 N37369 0 diode
R37370 N37369 N37370 10
D37370 N37370 0 diode
R37371 N37370 N37371 10
D37371 N37371 0 diode
R37372 N37371 N37372 10
D37372 N37372 0 diode
R37373 N37372 N37373 10
D37373 N37373 0 diode
R37374 N37373 N37374 10
D37374 N37374 0 diode
R37375 N37374 N37375 10
D37375 N37375 0 diode
R37376 N37375 N37376 10
D37376 N37376 0 diode
R37377 N37376 N37377 10
D37377 N37377 0 diode
R37378 N37377 N37378 10
D37378 N37378 0 diode
R37379 N37378 N37379 10
D37379 N37379 0 diode
R37380 N37379 N37380 10
D37380 N37380 0 diode
R37381 N37380 N37381 10
D37381 N37381 0 diode
R37382 N37381 N37382 10
D37382 N37382 0 diode
R37383 N37382 N37383 10
D37383 N37383 0 diode
R37384 N37383 N37384 10
D37384 N37384 0 diode
R37385 N37384 N37385 10
D37385 N37385 0 diode
R37386 N37385 N37386 10
D37386 N37386 0 diode
R37387 N37386 N37387 10
D37387 N37387 0 diode
R37388 N37387 N37388 10
D37388 N37388 0 diode
R37389 N37388 N37389 10
D37389 N37389 0 diode
R37390 N37389 N37390 10
D37390 N37390 0 diode
R37391 N37390 N37391 10
D37391 N37391 0 diode
R37392 N37391 N37392 10
D37392 N37392 0 diode
R37393 N37392 N37393 10
D37393 N37393 0 diode
R37394 N37393 N37394 10
D37394 N37394 0 diode
R37395 N37394 N37395 10
D37395 N37395 0 diode
R37396 N37395 N37396 10
D37396 N37396 0 diode
R37397 N37396 N37397 10
D37397 N37397 0 diode
R37398 N37397 N37398 10
D37398 N37398 0 diode
R37399 N37398 N37399 10
D37399 N37399 0 diode
R37400 N37399 N37400 10
D37400 N37400 0 diode
R37401 N37400 N37401 10
D37401 N37401 0 diode
R37402 N37401 N37402 10
D37402 N37402 0 diode
R37403 N37402 N37403 10
D37403 N37403 0 diode
R37404 N37403 N37404 10
D37404 N37404 0 diode
R37405 N37404 N37405 10
D37405 N37405 0 diode
R37406 N37405 N37406 10
D37406 N37406 0 diode
R37407 N37406 N37407 10
D37407 N37407 0 diode
R37408 N37407 N37408 10
D37408 N37408 0 diode
R37409 N37408 N37409 10
D37409 N37409 0 diode
R37410 N37409 N37410 10
D37410 N37410 0 diode
R37411 N37410 N37411 10
D37411 N37411 0 diode
R37412 N37411 N37412 10
D37412 N37412 0 diode
R37413 N37412 N37413 10
D37413 N37413 0 diode
R37414 N37413 N37414 10
D37414 N37414 0 diode
R37415 N37414 N37415 10
D37415 N37415 0 diode
R37416 N37415 N37416 10
D37416 N37416 0 diode
R37417 N37416 N37417 10
D37417 N37417 0 diode
R37418 N37417 N37418 10
D37418 N37418 0 diode
R37419 N37418 N37419 10
D37419 N37419 0 diode
R37420 N37419 N37420 10
D37420 N37420 0 diode
R37421 N37420 N37421 10
D37421 N37421 0 diode
R37422 N37421 N37422 10
D37422 N37422 0 diode
R37423 N37422 N37423 10
D37423 N37423 0 diode
R37424 N37423 N37424 10
D37424 N37424 0 diode
R37425 N37424 N37425 10
D37425 N37425 0 diode
R37426 N37425 N37426 10
D37426 N37426 0 diode
R37427 N37426 N37427 10
D37427 N37427 0 diode
R37428 N37427 N37428 10
D37428 N37428 0 diode
R37429 N37428 N37429 10
D37429 N37429 0 diode
R37430 N37429 N37430 10
D37430 N37430 0 diode
R37431 N37430 N37431 10
D37431 N37431 0 diode
R37432 N37431 N37432 10
D37432 N37432 0 diode
R37433 N37432 N37433 10
D37433 N37433 0 diode
R37434 N37433 N37434 10
D37434 N37434 0 diode
R37435 N37434 N37435 10
D37435 N37435 0 diode
R37436 N37435 N37436 10
D37436 N37436 0 diode
R37437 N37436 N37437 10
D37437 N37437 0 diode
R37438 N37437 N37438 10
D37438 N37438 0 diode
R37439 N37438 N37439 10
D37439 N37439 0 diode
R37440 N37439 N37440 10
D37440 N37440 0 diode
R37441 N37440 N37441 10
D37441 N37441 0 diode
R37442 N37441 N37442 10
D37442 N37442 0 diode
R37443 N37442 N37443 10
D37443 N37443 0 diode
R37444 N37443 N37444 10
D37444 N37444 0 diode
R37445 N37444 N37445 10
D37445 N37445 0 diode
R37446 N37445 N37446 10
D37446 N37446 0 diode
R37447 N37446 N37447 10
D37447 N37447 0 diode
R37448 N37447 N37448 10
D37448 N37448 0 diode
R37449 N37448 N37449 10
D37449 N37449 0 diode
R37450 N37449 N37450 10
D37450 N37450 0 diode
R37451 N37450 N37451 10
D37451 N37451 0 diode
R37452 N37451 N37452 10
D37452 N37452 0 diode
R37453 N37452 N37453 10
D37453 N37453 0 diode
R37454 N37453 N37454 10
D37454 N37454 0 diode
R37455 N37454 N37455 10
D37455 N37455 0 diode
R37456 N37455 N37456 10
D37456 N37456 0 diode
R37457 N37456 N37457 10
D37457 N37457 0 diode
R37458 N37457 N37458 10
D37458 N37458 0 diode
R37459 N37458 N37459 10
D37459 N37459 0 diode
R37460 N37459 N37460 10
D37460 N37460 0 diode
R37461 N37460 N37461 10
D37461 N37461 0 diode
R37462 N37461 N37462 10
D37462 N37462 0 diode
R37463 N37462 N37463 10
D37463 N37463 0 diode
R37464 N37463 N37464 10
D37464 N37464 0 diode
R37465 N37464 N37465 10
D37465 N37465 0 diode
R37466 N37465 N37466 10
D37466 N37466 0 diode
R37467 N37466 N37467 10
D37467 N37467 0 diode
R37468 N37467 N37468 10
D37468 N37468 0 diode
R37469 N37468 N37469 10
D37469 N37469 0 diode
R37470 N37469 N37470 10
D37470 N37470 0 diode
R37471 N37470 N37471 10
D37471 N37471 0 diode
R37472 N37471 N37472 10
D37472 N37472 0 diode
R37473 N37472 N37473 10
D37473 N37473 0 diode
R37474 N37473 N37474 10
D37474 N37474 0 diode
R37475 N37474 N37475 10
D37475 N37475 0 diode
R37476 N37475 N37476 10
D37476 N37476 0 diode
R37477 N37476 N37477 10
D37477 N37477 0 diode
R37478 N37477 N37478 10
D37478 N37478 0 diode
R37479 N37478 N37479 10
D37479 N37479 0 diode
R37480 N37479 N37480 10
D37480 N37480 0 diode
R37481 N37480 N37481 10
D37481 N37481 0 diode
R37482 N37481 N37482 10
D37482 N37482 0 diode
R37483 N37482 N37483 10
D37483 N37483 0 diode
R37484 N37483 N37484 10
D37484 N37484 0 diode
R37485 N37484 N37485 10
D37485 N37485 0 diode
R37486 N37485 N37486 10
D37486 N37486 0 diode
R37487 N37486 N37487 10
D37487 N37487 0 diode
R37488 N37487 N37488 10
D37488 N37488 0 diode
R37489 N37488 N37489 10
D37489 N37489 0 diode
R37490 N37489 N37490 10
D37490 N37490 0 diode
R37491 N37490 N37491 10
D37491 N37491 0 diode
R37492 N37491 N37492 10
D37492 N37492 0 diode
R37493 N37492 N37493 10
D37493 N37493 0 diode
R37494 N37493 N37494 10
D37494 N37494 0 diode
R37495 N37494 N37495 10
D37495 N37495 0 diode
R37496 N37495 N37496 10
D37496 N37496 0 diode
R37497 N37496 N37497 10
D37497 N37497 0 diode
R37498 N37497 N37498 10
D37498 N37498 0 diode
R37499 N37498 N37499 10
D37499 N37499 0 diode
R37500 N37499 N37500 10
D37500 N37500 0 diode
R37501 N37500 N37501 10
D37501 N37501 0 diode
R37502 N37501 N37502 10
D37502 N37502 0 diode
R37503 N37502 N37503 10
D37503 N37503 0 diode
R37504 N37503 N37504 10
D37504 N37504 0 diode
R37505 N37504 N37505 10
D37505 N37505 0 diode
R37506 N37505 N37506 10
D37506 N37506 0 diode
R37507 N37506 N37507 10
D37507 N37507 0 diode
R37508 N37507 N37508 10
D37508 N37508 0 diode
R37509 N37508 N37509 10
D37509 N37509 0 diode
R37510 N37509 N37510 10
D37510 N37510 0 diode
R37511 N37510 N37511 10
D37511 N37511 0 diode
R37512 N37511 N37512 10
D37512 N37512 0 diode
R37513 N37512 N37513 10
D37513 N37513 0 diode
R37514 N37513 N37514 10
D37514 N37514 0 diode
R37515 N37514 N37515 10
D37515 N37515 0 diode
R37516 N37515 N37516 10
D37516 N37516 0 diode
R37517 N37516 N37517 10
D37517 N37517 0 diode
R37518 N37517 N37518 10
D37518 N37518 0 diode
R37519 N37518 N37519 10
D37519 N37519 0 diode
R37520 N37519 N37520 10
D37520 N37520 0 diode
R37521 N37520 N37521 10
D37521 N37521 0 diode
R37522 N37521 N37522 10
D37522 N37522 0 diode
R37523 N37522 N37523 10
D37523 N37523 0 diode
R37524 N37523 N37524 10
D37524 N37524 0 diode
R37525 N37524 N37525 10
D37525 N37525 0 diode
R37526 N37525 N37526 10
D37526 N37526 0 diode
R37527 N37526 N37527 10
D37527 N37527 0 diode
R37528 N37527 N37528 10
D37528 N37528 0 diode
R37529 N37528 N37529 10
D37529 N37529 0 diode
R37530 N37529 N37530 10
D37530 N37530 0 diode
R37531 N37530 N37531 10
D37531 N37531 0 diode
R37532 N37531 N37532 10
D37532 N37532 0 diode
R37533 N37532 N37533 10
D37533 N37533 0 diode
R37534 N37533 N37534 10
D37534 N37534 0 diode
R37535 N37534 N37535 10
D37535 N37535 0 diode
R37536 N37535 N37536 10
D37536 N37536 0 diode
R37537 N37536 N37537 10
D37537 N37537 0 diode
R37538 N37537 N37538 10
D37538 N37538 0 diode
R37539 N37538 N37539 10
D37539 N37539 0 diode
R37540 N37539 N37540 10
D37540 N37540 0 diode
R37541 N37540 N37541 10
D37541 N37541 0 diode
R37542 N37541 N37542 10
D37542 N37542 0 diode
R37543 N37542 N37543 10
D37543 N37543 0 diode
R37544 N37543 N37544 10
D37544 N37544 0 diode
R37545 N37544 N37545 10
D37545 N37545 0 diode
R37546 N37545 N37546 10
D37546 N37546 0 diode
R37547 N37546 N37547 10
D37547 N37547 0 diode
R37548 N37547 N37548 10
D37548 N37548 0 diode
R37549 N37548 N37549 10
D37549 N37549 0 diode
R37550 N37549 N37550 10
D37550 N37550 0 diode
R37551 N37550 N37551 10
D37551 N37551 0 diode
R37552 N37551 N37552 10
D37552 N37552 0 diode
R37553 N37552 N37553 10
D37553 N37553 0 diode
R37554 N37553 N37554 10
D37554 N37554 0 diode
R37555 N37554 N37555 10
D37555 N37555 0 diode
R37556 N37555 N37556 10
D37556 N37556 0 diode
R37557 N37556 N37557 10
D37557 N37557 0 diode
R37558 N37557 N37558 10
D37558 N37558 0 diode
R37559 N37558 N37559 10
D37559 N37559 0 diode
R37560 N37559 N37560 10
D37560 N37560 0 diode
R37561 N37560 N37561 10
D37561 N37561 0 diode
R37562 N37561 N37562 10
D37562 N37562 0 diode
R37563 N37562 N37563 10
D37563 N37563 0 diode
R37564 N37563 N37564 10
D37564 N37564 0 diode
R37565 N37564 N37565 10
D37565 N37565 0 diode
R37566 N37565 N37566 10
D37566 N37566 0 diode
R37567 N37566 N37567 10
D37567 N37567 0 diode
R37568 N37567 N37568 10
D37568 N37568 0 diode
R37569 N37568 N37569 10
D37569 N37569 0 diode
R37570 N37569 N37570 10
D37570 N37570 0 diode
R37571 N37570 N37571 10
D37571 N37571 0 diode
R37572 N37571 N37572 10
D37572 N37572 0 diode
R37573 N37572 N37573 10
D37573 N37573 0 diode
R37574 N37573 N37574 10
D37574 N37574 0 diode
R37575 N37574 N37575 10
D37575 N37575 0 diode
R37576 N37575 N37576 10
D37576 N37576 0 diode
R37577 N37576 N37577 10
D37577 N37577 0 diode
R37578 N37577 N37578 10
D37578 N37578 0 diode
R37579 N37578 N37579 10
D37579 N37579 0 diode
R37580 N37579 N37580 10
D37580 N37580 0 diode
R37581 N37580 N37581 10
D37581 N37581 0 diode
R37582 N37581 N37582 10
D37582 N37582 0 diode
R37583 N37582 N37583 10
D37583 N37583 0 diode
R37584 N37583 N37584 10
D37584 N37584 0 diode
R37585 N37584 N37585 10
D37585 N37585 0 diode
R37586 N37585 N37586 10
D37586 N37586 0 diode
R37587 N37586 N37587 10
D37587 N37587 0 diode
R37588 N37587 N37588 10
D37588 N37588 0 diode
R37589 N37588 N37589 10
D37589 N37589 0 diode
R37590 N37589 N37590 10
D37590 N37590 0 diode
R37591 N37590 N37591 10
D37591 N37591 0 diode
R37592 N37591 N37592 10
D37592 N37592 0 diode
R37593 N37592 N37593 10
D37593 N37593 0 diode
R37594 N37593 N37594 10
D37594 N37594 0 diode
R37595 N37594 N37595 10
D37595 N37595 0 diode
R37596 N37595 N37596 10
D37596 N37596 0 diode
R37597 N37596 N37597 10
D37597 N37597 0 diode
R37598 N37597 N37598 10
D37598 N37598 0 diode
R37599 N37598 N37599 10
D37599 N37599 0 diode
R37600 N37599 N37600 10
D37600 N37600 0 diode
R37601 N37600 N37601 10
D37601 N37601 0 diode
R37602 N37601 N37602 10
D37602 N37602 0 diode
R37603 N37602 N37603 10
D37603 N37603 0 diode
R37604 N37603 N37604 10
D37604 N37604 0 diode
R37605 N37604 N37605 10
D37605 N37605 0 diode
R37606 N37605 N37606 10
D37606 N37606 0 diode
R37607 N37606 N37607 10
D37607 N37607 0 diode
R37608 N37607 N37608 10
D37608 N37608 0 diode
R37609 N37608 N37609 10
D37609 N37609 0 diode
R37610 N37609 N37610 10
D37610 N37610 0 diode
R37611 N37610 N37611 10
D37611 N37611 0 diode
R37612 N37611 N37612 10
D37612 N37612 0 diode
R37613 N37612 N37613 10
D37613 N37613 0 diode
R37614 N37613 N37614 10
D37614 N37614 0 diode
R37615 N37614 N37615 10
D37615 N37615 0 diode
R37616 N37615 N37616 10
D37616 N37616 0 diode
R37617 N37616 N37617 10
D37617 N37617 0 diode
R37618 N37617 N37618 10
D37618 N37618 0 diode
R37619 N37618 N37619 10
D37619 N37619 0 diode
R37620 N37619 N37620 10
D37620 N37620 0 diode
R37621 N37620 N37621 10
D37621 N37621 0 diode
R37622 N37621 N37622 10
D37622 N37622 0 diode
R37623 N37622 N37623 10
D37623 N37623 0 diode
R37624 N37623 N37624 10
D37624 N37624 0 diode
R37625 N37624 N37625 10
D37625 N37625 0 diode
R37626 N37625 N37626 10
D37626 N37626 0 diode
R37627 N37626 N37627 10
D37627 N37627 0 diode
R37628 N37627 N37628 10
D37628 N37628 0 diode
R37629 N37628 N37629 10
D37629 N37629 0 diode
R37630 N37629 N37630 10
D37630 N37630 0 diode
R37631 N37630 N37631 10
D37631 N37631 0 diode
R37632 N37631 N37632 10
D37632 N37632 0 diode
R37633 N37632 N37633 10
D37633 N37633 0 diode
R37634 N37633 N37634 10
D37634 N37634 0 diode
R37635 N37634 N37635 10
D37635 N37635 0 diode
R37636 N37635 N37636 10
D37636 N37636 0 diode
R37637 N37636 N37637 10
D37637 N37637 0 diode
R37638 N37637 N37638 10
D37638 N37638 0 diode
R37639 N37638 N37639 10
D37639 N37639 0 diode
R37640 N37639 N37640 10
D37640 N37640 0 diode
R37641 N37640 N37641 10
D37641 N37641 0 diode
R37642 N37641 N37642 10
D37642 N37642 0 diode
R37643 N37642 N37643 10
D37643 N37643 0 diode
R37644 N37643 N37644 10
D37644 N37644 0 diode
R37645 N37644 N37645 10
D37645 N37645 0 diode
R37646 N37645 N37646 10
D37646 N37646 0 diode
R37647 N37646 N37647 10
D37647 N37647 0 diode
R37648 N37647 N37648 10
D37648 N37648 0 diode
R37649 N37648 N37649 10
D37649 N37649 0 diode
R37650 N37649 N37650 10
D37650 N37650 0 diode
R37651 N37650 N37651 10
D37651 N37651 0 diode
R37652 N37651 N37652 10
D37652 N37652 0 diode
R37653 N37652 N37653 10
D37653 N37653 0 diode
R37654 N37653 N37654 10
D37654 N37654 0 diode
R37655 N37654 N37655 10
D37655 N37655 0 diode
R37656 N37655 N37656 10
D37656 N37656 0 diode
R37657 N37656 N37657 10
D37657 N37657 0 diode
R37658 N37657 N37658 10
D37658 N37658 0 diode
R37659 N37658 N37659 10
D37659 N37659 0 diode
R37660 N37659 N37660 10
D37660 N37660 0 diode
R37661 N37660 N37661 10
D37661 N37661 0 diode
R37662 N37661 N37662 10
D37662 N37662 0 diode
R37663 N37662 N37663 10
D37663 N37663 0 diode
R37664 N37663 N37664 10
D37664 N37664 0 diode
R37665 N37664 N37665 10
D37665 N37665 0 diode
R37666 N37665 N37666 10
D37666 N37666 0 diode
R37667 N37666 N37667 10
D37667 N37667 0 diode
R37668 N37667 N37668 10
D37668 N37668 0 diode
R37669 N37668 N37669 10
D37669 N37669 0 diode
R37670 N37669 N37670 10
D37670 N37670 0 diode
R37671 N37670 N37671 10
D37671 N37671 0 diode
R37672 N37671 N37672 10
D37672 N37672 0 diode
R37673 N37672 N37673 10
D37673 N37673 0 diode
R37674 N37673 N37674 10
D37674 N37674 0 diode
R37675 N37674 N37675 10
D37675 N37675 0 diode
R37676 N37675 N37676 10
D37676 N37676 0 diode
R37677 N37676 N37677 10
D37677 N37677 0 diode
R37678 N37677 N37678 10
D37678 N37678 0 diode
R37679 N37678 N37679 10
D37679 N37679 0 diode
R37680 N37679 N37680 10
D37680 N37680 0 diode
R37681 N37680 N37681 10
D37681 N37681 0 diode
R37682 N37681 N37682 10
D37682 N37682 0 diode
R37683 N37682 N37683 10
D37683 N37683 0 diode
R37684 N37683 N37684 10
D37684 N37684 0 diode
R37685 N37684 N37685 10
D37685 N37685 0 diode
R37686 N37685 N37686 10
D37686 N37686 0 diode
R37687 N37686 N37687 10
D37687 N37687 0 diode
R37688 N37687 N37688 10
D37688 N37688 0 diode
R37689 N37688 N37689 10
D37689 N37689 0 diode
R37690 N37689 N37690 10
D37690 N37690 0 diode
R37691 N37690 N37691 10
D37691 N37691 0 diode
R37692 N37691 N37692 10
D37692 N37692 0 diode
R37693 N37692 N37693 10
D37693 N37693 0 diode
R37694 N37693 N37694 10
D37694 N37694 0 diode
R37695 N37694 N37695 10
D37695 N37695 0 diode
R37696 N37695 N37696 10
D37696 N37696 0 diode
R37697 N37696 N37697 10
D37697 N37697 0 diode
R37698 N37697 N37698 10
D37698 N37698 0 diode
R37699 N37698 N37699 10
D37699 N37699 0 diode
R37700 N37699 N37700 10
D37700 N37700 0 diode
R37701 N37700 N37701 10
D37701 N37701 0 diode
R37702 N37701 N37702 10
D37702 N37702 0 diode
R37703 N37702 N37703 10
D37703 N37703 0 diode
R37704 N37703 N37704 10
D37704 N37704 0 diode
R37705 N37704 N37705 10
D37705 N37705 0 diode
R37706 N37705 N37706 10
D37706 N37706 0 diode
R37707 N37706 N37707 10
D37707 N37707 0 diode
R37708 N37707 N37708 10
D37708 N37708 0 diode
R37709 N37708 N37709 10
D37709 N37709 0 diode
R37710 N37709 N37710 10
D37710 N37710 0 diode
R37711 N37710 N37711 10
D37711 N37711 0 diode
R37712 N37711 N37712 10
D37712 N37712 0 diode
R37713 N37712 N37713 10
D37713 N37713 0 diode
R37714 N37713 N37714 10
D37714 N37714 0 diode
R37715 N37714 N37715 10
D37715 N37715 0 diode
R37716 N37715 N37716 10
D37716 N37716 0 diode
R37717 N37716 N37717 10
D37717 N37717 0 diode
R37718 N37717 N37718 10
D37718 N37718 0 diode
R37719 N37718 N37719 10
D37719 N37719 0 diode
R37720 N37719 N37720 10
D37720 N37720 0 diode
R37721 N37720 N37721 10
D37721 N37721 0 diode
R37722 N37721 N37722 10
D37722 N37722 0 diode
R37723 N37722 N37723 10
D37723 N37723 0 diode
R37724 N37723 N37724 10
D37724 N37724 0 diode
R37725 N37724 N37725 10
D37725 N37725 0 diode
R37726 N37725 N37726 10
D37726 N37726 0 diode
R37727 N37726 N37727 10
D37727 N37727 0 diode
R37728 N37727 N37728 10
D37728 N37728 0 diode
R37729 N37728 N37729 10
D37729 N37729 0 diode
R37730 N37729 N37730 10
D37730 N37730 0 diode
R37731 N37730 N37731 10
D37731 N37731 0 diode
R37732 N37731 N37732 10
D37732 N37732 0 diode
R37733 N37732 N37733 10
D37733 N37733 0 diode
R37734 N37733 N37734 10
D37734 N37734 0 diode
R37735 N37734 N37735 10
D37735 N37735 0 diode
R37736 N37735 N37736 10
D37736 N37736 0 diode
R37737 N37736 N37737 10
D37737 N37737 0 diode
R37738 N37737 N37738 10
D37738 N37738 0 diode
R37739 N37738 N37739 10
D37739 N37739 0 diode
R37740 N37739 N37740 10
D37740 N37740 0 diode
R37741 N37740 N37741 10
D37741 N37741 0 diode
R37742 N37741 N37742 10
D37742 N37742 0 diode
R37743 N37742 N37743 10
D37743 N37743 0 diode
R37744 N37743 N37744 10
D37744 N37744 0 diode
R37745 N37744 N37745 10
D37745 N37745 0 diode
R37746 N37745 N37746 10
D37746 N37746 0 diode
R37747 N37746 N37747 10
D37747 N37747 0 diode
R37748 N37747 N37748 10
D37748 N37748 0 diode
R37749 N37748 N37749 10
D37749 N37749 0 diode
R37750 N37749 N37750 10
D37750 N37750 0 diode
R37751 N37750 N37751 10
D37751 N37751 0 diode
R37752 N37751 N37752 10
D37752 N37752 0 diode
R37753 N37752 N37753 10
D37753 N37753 0 diode
R37754 N37753 N37754 10
D37754 N37754 0 diode
R37755 N37754 N37755 10
D37755 N37755 0 diode
R37756 N37755 N37756 10
D37756 N37756 0 diode
R37757 N37756 N37757 10
D37757 N37757 0 diode
R37758 N37757 N37758 10
D37758 N37758 0 diode
R37759 N37758 N37759 10
D37759 N37759 0 diode
R37760 N37759 N37760 10
D37760 N37760 0 diode
R37761 N37760 N37761 10
D37761 N37761 0 diode
R37762 N37761 N37762 10
D37762 N37762 0 diode
R37763 N37762 N37763 10
D37763 N37763 0 diode
R37764 N37763 N37764 10
D37764 N37764 0 diode
R37765 N37764 N37765 10
D37765 N37765 0 diode
R37766 N37765 N37766 10
D37766 N37766 0 diode
R37767 N37766 N37767 10
D37767 N37767 0 diode
R37768 N37767 N37768 10
D37768 N37768 0 diode
R37769 N37768 N37769 10
D37769 N37769 0 diode
R37770 N37769 N37770 10
D37770 N37770 0 diode
R37771 N37770 N37771 10
D37771 N37771 0 diode
R37772 N37771 N37772 10
D37772 N37772 0 diode
R37773 N37772 N37773 10
D37773 N37773 0 diode
R37774 N37773 N37774 10
D37774 N37774 0 diode
R37775 N37774 N37775 10
D37775 N37775 0 diode
R37776 N37775 N37776 10
D37776 N37776 0 diode
R37777 N37776 N37777 10
D37777 N37777 0 diode
R37778 N37777 N37778 10
D37778 N37778 0 diode
R37779 N37778 N37779 10
D37779 N37779 0 diode
R37780 N37779 N37780 10
D37780 N37780 0 diode
R37781 N37780 N37781 10
D37781 N37781 0 diode
R37782 N37781 N37782 10
D37782 N37782 0 diode
R37783 N37782 N37783 10
D37783 N37783 0 diode
R37784 N37783 N37784 10
D37784 N37784 0 diode
R37785 N37784 N37785 10
D37785 N37785 0 diode
R37786 N37785 N37786 10
D37786 N37786 0 diode
R37787 N37786 N37787 10
D37787 N37787 0 diode
R37788 N37787 N37788 10
D37788 N37788 0 diode
R37789 N37788 N37789 10
D37789 N37789 0 diode
R37790 N37789 N37790 10
D37790 N37790 0 diode
R37791 N37790 N37791 10
D37791 N37791 0 diode
R37792 N37791 N37792 10
D37792 N37792 0 diode
R37793 N37792 N37793 10
D37793 N37793 0 diode
R37794 N37793 N37794 10
D37794 N37794 0 diode
R37795 N37794 N37795 10
D37795 N37795 0 diode
R37796 N37795 N37796 10
D37796 N37796 0 diode
R37797 N37796 N37797 10
D37797 N37797 0 diode
R37798 N37797 N37798 10
D37798 N37798 0 diode
R37799 N37798 N37799 10
D37799 N37799 0 diode
R37800 N37799 N37800 10
D37800 N37800 0 diode
R37801 N37800 N37801 10
D37801 N37801 0 diode
R37802 N37801 N37802 10
D37802 N37802 0 diode
R37803 N37802 N37803 10
D37803 N37803 0 diode
R37804 N37803 N37804 10
D37804 N37804 0 diode
R37805 N37804 N37805 10
D37805 N37805 0 diode
R37806 N37805 N37806 10
D37806 N37806 0 diode
R37807 N37806 N37807 10
D37807 N37807 0 diode
R37808 N37807 N37808 10
D37808 N37808 0 diode
R37809 N37808 N37809 10
D37809 N37809 0 diode
R37810 N37809 N37810 10
D37810 N37810 0 diode
R37811 N37810 N37811 10
D37811 N37811 0 diode
R37812 N37811 N37812 10
D37812 N37812 0 diode
R37813 N37812 N37813 10
D37813 N37813 0 diode
R37814 N37813 N37814 10
D37814 N37814 0 diode
R37815 N37814 N37815 10
D37815 N37815 0 diode
R37816 N37815 N37816 10
D37816 N37816 0 diode
R37817 N37816 N37817 10
D37817 N37817 0 diode
R37818 N37817 N37818 10
D37818 N37818 0 diode
R37819 N37818 N37819 10
D37819 N37819 0 diode
R37820 N37819 N37820 10
D37820 N37820 0 diode
R37821 N37820 N37821 10
D37821 N37821 0 diode
R37822 N37821 N37822 10
D37822 N37822 0 diode
R37823 N37822 N37823 10
D37823 N37823 0 diode
R37824 N37823 N37824 10
D37824 N37824 0 diode
R37825 N37824 N37825 10
D37825 N37825 0 diode
R37826 N37825 N37826 10
D37826 N37826 0 diode
R37827 N37826 N37827 10
D37827 N37827 0 diode
R37828 N37827 N37828 10
D37828 N37828 0 diode
R37829 N37828 N37829 10
D37829 N37829 0 diode
R37830 N37829 N37830 10
D37830 N37830 0 diode
R37831 N37830 N37831 10
D37831 N37831 0 diode
R37832 N37831 N37832 10
D37832 N37832 0 diode
R37833 N37832 N37833 10
D37833 N37833 0 diode
R37834 N37833 N37834 10
D37834 N37834 0 diode
R37835 N37834 N37835 10
D37835 N37835 0 diode
R37836 N37835 N37836 10
D37836 N37836 0 diode
R37837 N37836 N37837 10
D37837 N37837 0 diode
R37838 N37837 N37838 10
D37838 N37838 0 diode
R37839 N37838 N37839 10
D37839 N37839 0 diode
R37840 N37839 N37840 10
D37840 N37840 0 diode
R37841 N37840 N37841 10
D37841 N37841 0 diode
R37842 N37841 N37842 10
D37842 N37842 0 diode
R37843 N37842 N37843 10
D37843 N37843 0 diode
R37844 N37843 N37844 10
D37844 N37844 0 diode
R37845 N37844 N37845 10
D37845 N37845 0 diode
R37846 N37845 N37846 10
D37846 N37846 0 diode
R37847 N37846 N37847 10
D37847 N37847 0 diode
R37848 N37847 N37848 10
D37848 N37848 0 diode
R37849 N37848 N37849 10
D37849 N37849 0 diode
R37850 N37849 N37850 10
D37850 N37850 0 diode
R37851 N37850 N37851 10
D37851 N37851 0 diode
R37852 N37851 N37852 10
D37852 N37852 0 diode
R37853 N37852 N37853 10
D37853 N37853 0 diode
R37854 N37853 N37854 10
D37854 N37854 0 diode
R37855 N37854 N37855 10
D37855 N37855 0 diode
R37856 N37855 N37856 10
D37856 N37856 0 diode
R37857 N37856 N37857 10
D37857 N37857 0 diode
R37858 N37857 N37858 10
D37858 N37858 0 diode
R37859 N37858 N37859 10
D37859 N37859 0 diode
R37860 N37859 N37860 10
D37860 N37860 0 diode
R37861 N37860 N37861 10
D37861 N37861 0 diode
R37862 N37861 N37862 10
D37862 N37862 0 diode
R37863 N37862 N37863 10
D37863 N37863 0 diode
R37864 N37863 N37864 10
D37864 N37864 0 diode
R37865 N37864 N37865 10
D37865 N37865 0 diode
R37866 N37865 N37866 10
D37866 N37866 0 diode
R37867 N37866 N37867 10
D37867 N37867 0 diode
R37868 N37867 N37868 10
D37868 N37868 0 diode
R37869 N37868 N37869 10
D37869 N37869 0 diode
R37870 N37869 N37870 10
D37870 N37870 0 diode
R37871 N37870 N37871 10
D37871 N37871 0 diode
R37872 N37871 N37872 10
D37872 N37872 0 diode
R37873 N37872 N37873 10
D37873 N37873 0 diode
R37874 N37873 N37874 10
D37874 N37874 0 diode
R37875 N37874 N37875 10
D37875 N37875 0 diode
R37876 N37875 N37876 10
D37876 N37876 0 diode
R37877 N37876 N37877 10
D37877 N37877 0 diode
R37878 N37877 N37878 10
D37878 N37878 0 diode
R37879 N37878 N37879 10
D37879 N37879 0 diode
R37880 N37879 N37880 10
D37880 N37880 0 diode
R37881 N37880 N37881 10
D37881 N37881 0 diode
R37882 N37881 N37882 10
D37882 N37882 0 diode
R37883 N37882 N37883 10
D37883 N37883 0 diode
R37884 N37883 N37884 10
D37884 N37884 0 diode
R37885 N37884 N37885 10
D37885 N37885 0 diode
R37886 N37885 N37886 10
D37886 N37886 0 diode
R37887 N37886 N37887 10
D37887 N37887 0 diode
R37888 N37887 N37888 10
D37888 N37888 0 diode
R37889 N37888 N37889 10
D37889 N37889 0 diode
R37890 N37889 N37890 10
D37890 N37890 0 diode
R37891 N37890 N37891 10
D37891 N37891 0 diode
R37892 N37891 N37892 10
D37892 N37892 0 diode
R37893 N37892 N37893 10
D37893 N37893 0 diode
R37894 N37893 N37894 10
D37894 N37894 0 diode
R37895 N37894 N37895 10
D37895 N37895 0 diode
R37896 N37895 N37896 10
D37896 N37896 0 diode
R37897 N37896 N37897 10
D37897 N37897 0 diode
R37898 N37897 N37898 10
D37898 N37898 0 diode
R37899 N37898 N37899 10
D37899 N37899 0 diode
R37900 N37899 N37900 10
D37900 N37900 0 diode
R37901 N37900 N37901 10
D37901 N37901 0 diode
R37902 N37901 N37902 10
D37902 N37902 0 diode
R37903 N37902 N37903 10
D37903 N37903 0 diode
R37904 N37903 N37904 10
D37904 N37904 0 diode
R37905 N37904 N37905 10
D37905 N37905 0 diode
R37906 N37905 N37906 10
D37906 N37906 0 diode
R37907 N37906 N37907 10
D37907 N37907 0 diode
R37908 N37907 N37908 10
D37908 N37908 0 diode
R37909 N37908 N37909 10
D37909 N37909 0 diode
R37910 N37909 N37910 10
D37910 N37910 0 diode
R37911 N37910 N37911 10
D37911 N37911 0 diode
R37912 N37911 N37912 10
D37912 N37912 0 diode
R37913 N37912 N37913 10
D37913 N37913 0 diode
R37914 N37913 N37914 10
D37914 N37914 0 diode
R37915 N37914 N37915 10
D37915 N37915 0 diode
R37916 N37915 N37916 10
D37916 N37916 0 diode
R37917 N37916 N37917 10
D37917 N37917 0 diode
R37918 N37917 N37918 10
D37918 N37918 0 diode
R37919 N37918 N37919 10
D37919 N37919 0 diode
R37920 N37919 N37920 10
D37920 N37920 0 diode
R37921 N37920 N37921 10
D37921 N37921 0 diode
R37922 N37921 N37922 10
D37922 N37922 0 diode
R37923 N37922 N37923 10
D37923 N37923 0 diode
R37924 N37923 N37924 10
D37924 N37924 0 diode
R37925 N37924 N37925 10
D37925 N37925 0 diode
R37926 N37925 N37926 10
D37926 N37926 0 diode
R37927 N37926 N37927 10
D37927 N37927 0 diode
R37928 N37927 N37928 10
D37928 N37928 0 diode
R37929 N37928 N37929 10
D37929 N37929 0 diode
R37930 N37929 N37930 10
D37930 N37930 0 diode
R37931 N37930 N37931 10
D37931 N37931 0 diode
R37932 N37931 N37932 10
D37932 N37932 0 diode
R37933 N37932 N37933 10
D37933 N37933 0 diode
R37934 N37933 N37934 10
D37934 N37934 0 diode
R37935 N37934 N37935 10
D37935 N37935 0 diode
R37936 N37935 N37936 10
D37936 N37936 0 diode
R37937 N37936 N37937 10
D37937 N37937 0 diode
R37938 N37937 N37938 10
D37938 N37938 0 diode
R37939 N37938 N37939 10
D37939 N37939 0 diode
R37940 N37939 N37940 10
D37940 N37940 0 diode
R37941 N37940 N37941 10
D37941 N37941 0 diode
R37942 N37941 N37942 10
D37942 N37942 0 diode
R37943 N37942 N37943 10
D37943 N37943 0 diode
R37944 N37943 N37944 10
D37944 N37944 0 diode
R37945 N37944 N37945 10
D37945 N37945 0 diode
R37946 N37945 N37946 10
D37946 N37946 0 diode
R37947 N37946 N37947 10
D37947 N37947 0 diode
R37948 N37947 N37948 10
D37948 N37948 0 diode
R37949 N37948 N37949 10
D37949 N37949 0 diode
R37950 N37949 N37950 10
D37950 N37950 0 diode
R37951 N37950 N37951 10
D37951 N37951 0 diode
R37952 N37951 N37952 10
D37952 N37952 0 diode
R37953 N37952 N37953 10
D37953 N37953 0 diode
R37954 N37953 N37954 10
D37954 N37954 0 diode
R37955 N37954 N37955 10
D37955 N37955 0 diode
R37956 N37955 N37956 10
D37956 N37956 0 diode
R37957 N37956 N37957 10
D37957 N37957 0 diode
R37958 N37957 N37958 10
D37958 N37958 0 diode
R37959 N37958 N37959 10
D37959 N37959 0 diode
R37960 N37959 N37960 10
D37960 N37960 0 diode
R37961 N37960 N37961 10
D37961 N37961 0 diode
R37962 N37961 N37962 10
D37962 N37962 0 diode
R37963 N37962 N37963 10
D37963 N37963 0 diode
R37964 N37963 N37964 10
D37964 N37964 0 diode
R37965 N37964 N37965 10
D37965 N37965 0 diode
R37966 N37965 N37966 10
D37966 N37966 0 diode
R37967 N37966 N37967 10
D37967 N37967 0 diode
R37968 N37967 N37968 10
D37968 N37968 0 diode
R37969 N37968 N37969 10
D37969 N37969 0 diode
R37970 N37969 N37970 10
D37970 N37970 0 diode
R37971 N37970 N37971 10
D37971 N37971 0 diode
R37972 N37971 N37972 10
D37972 N37972 0 diode
R37973 N37972 N37973 10
D37973 N37973 0 diode
R37974 N37973 N37974 10
D37974 N37974 0 diode
R37975 N37974 N37975 10
D37975 N37975 0 diode
R37976 N37975 N37976 10
D37976 N37976 0 diode
R37977 N37976 N37977 10
D37977 N37977 0 diode
R37978 N37977 N37978 10
D37978 N37978 0 diode
R37979 N37978 N37979 10
D37979 N37979 0 diode
R37980 N37979 N37980 10
D37980 N37980 0 diode
R37981 N37980 N37981 10
D37981 N37981 0 diode
R37982 N37981 N37982 10
D37982 N37982 0 diode
R37983 N37982 N37983 10
D37983 N37983 0 diode
R37984 N37983 N37984 10
D37984 N37984 0 diode
R37985 N37984 N37985 10
D37985 N37985 0 diode
R37986 N37985 N37986 10
D37986 N37986 0 diode
R37987 N37986 N37987 10
D37987 N37987 0 diode
R37988 N37987 N37988 10
D37988 N37988 0 diode
R37989 N37988 N37989 10
D37989 N37989 0 diode
R37990 N37989 N37990 10
D37990 N37990 0 diode
R37991 N37990 N37991 10
D37991 N37991 0 diode
R37992 N37991 N37992 10
D37992 N37992 0 diode
R37993 N37992 N37993 10
D37993 N37993 0 diode
R37994 N37993 N37994 10
D37994 N37994 0 diode
R37995 N37994 N37995 10
D37995 N37995 0 diode
R37996 N37995 N37996 10
D37996 N37996 0 diode
R37997 N37996 N37997 10
D37997 N37997 0 diode
R37998 N37997 N37998 10
D37998 N37998 0 diode
R37999 N37998 N37999 10
D37999 N37999 0 diode
R38000 N37999 N38000 10
D38000 N38000 0 diode
R38001 N38000 N38001 10
D38001 N38001 0 diode
R38002 N38001 N38002 10
D38002 N38002 0 diode
R38003 N38002 N38003 10
D38003 N38003 0 diode
R38004 N38003 N38004 10
D38004 N38004 0 diode
R38005 N38004 N38005 10
D38005 N38005 0 diode
R38006 N38005 N38006 10
D38006 N38006 0 diode
R38007 N38006 N38007 10
D38007 N38007 0 diode
R38008 N38007 N38008 10
D38008 N38008 0 diode
R38009 N38008 N38009 10
D38009 N38009 0 diode
R38010 N38009 N38010 10
D38010 N38010 0 diode
R38011 N38010 N38011 10
D38011 N38011 0 diode
R38012 N38011 N38012 10
D38012 N38012 0 diode
R38013 N38012 N38013 10
D38013 N38013 0 diode
R38014 N38013 N38014 10
D38014 N38014 0 diode
R38015 N38014 N38015 10
D38015 N38015 0 diode
R38016 N38015 N38016 10
D38016 N38016 0 diode
R38017 N38016 N38017 10
D38017 N38017 0 diode
R38018 N38017 N38018 10
D38018 N38018 0 diode
R38019 N38018 N38019 10
D38019 N38019 0 diode
R38020 N38019 N38020 10
D38020 N38020 0 diode
R38021 N38020 N38021 10
D38021 N38021 0 diode
R38022 N38021 N38022 10
D38022 N38022 0 diode
R38023 N38022 N38023 10
D38023 N38023 0 diode
R38024 N38023 N38024 10
D38024 N38024 0 diode
R38025 N38024 N38025 10
D38025 N38025 0 diode
R38026 N38025 N38026 10
D38026 N38026 0 diode
R38027 N38026 N38027 10
D38027 N38027 0 diode
R38028 N38027 N38028 10
D38028 N38028 0 diode
R38029 N38028 N38029 10
D38029 N38029 0 diode
R38030 N38029 N38030 10
D38030 N38030 0 diode
R38031 N38030 N38031 10
D38031 N38031 0 diode
R38032 N38031 N38032 10
D38032 N38032 0 diode
R38033 N38032 N38033 10
D38033 N38033 0 diode
R38034 N38033 N38034 10
D38034 N38034 0 diode
R38035 N38034 N38035 10
D38035 N38035 0 diode
R38036 N38035 N38036 10
D38036 N38036 0 diode
R38037 N38036 N38037 10
D38037 N38037 0 diode
R38038 N38037 N38038 10
D38038 N38038 0 diode
R38039 N38038 N38039 10
D38039 N38039 0 diode
R38040 N38039 N38040 10
D38040 N38040 0 diode
R38041 N38040 N38041 10
D38041 N38041 0 diode
R38042 N38041 N38042 10
D38042 N38042 0 diode
R38043 N38042 N38043 10
D38043 N38043 0 diode
R38044 N38043 N38044 10
D38044 N38044 0 diode
R38045 N38044 N38045 10
D38045 N38045 0 diode
R38046 N38045 N38046 10
D38046 N38046 0 diode
R38047 N38046 N38047 10
D38047 N38047 0 diode
R38048 N38047 N38048 10
D38048 N38048 0 diode
R38049 N38048 N38049 10
D38049 N38049 0 diode
R38050 N38049 N38050 10
D38050 N38050 0 diode
R38051 N38050 N38051 10
D38051 N38051 0 diode
R38052 N38051 N38052 10
D38052 N38052 0 diode
R38053 N38052 N38053 10
D38053 N38053 0 diode
R38054 N38053 N38054 10
D38054 N38054 0 diode
R38055 N38054 N38055 10
D38055 N38055 0 diode
R38056 N38055 N38056 10
D38056 N38056 0 diode
R38057 N38056 N38057 10
D38057 N38057 0 diode
R38058 N38057 N38058 10
D38058 N38058 0 diode
R38059 N38058 N38059 10
D38059 N38059 0 diode
R38060 N38059 N38060 10
D38060 N38060 0 diode
R38061 N38060 N38061 10
D38061 N38061 0 diode
R38062 N38061 N38062 10
D38062 N38062 0 diode
R38063 N38062 N38063 10
D38063 N38063 0 diode
R38064 N38063 N38064 10
D38064 N38064 0 diode
R38065 N38064 N38065 10
D38065 N38065 0 diode
R38066 N38065 N38066 10
D38066 N38066 0 diode
R38067 N38066 N38067 10
D38067 N38067 0 diode
R38068 N38067 N38068 10
D38068 N38068 0 diode
R38069 N38068 N38069 10
D38069 N38069 0 diode
R38070 N38069 N38070 10
D38070 N38070 0 diode
R38071 N38070 N38071 10
D38071 N38071 0 diode
R38072 N38071 N38072 10
D38072 N38072 0 diode
R38073 N38072 N38073 10
D38073 N38073 0 diode
R38074 N38073 N38074 10
D38074 N38074 0 diode
R38075 N38074 N38075 10
D38075 N38075 0 diode
R38076 N38075 N38076 10
D38076 N38076 0 diode
R38077 N38076 N38077 10
D38077 N38077 0 diode
R38078 N38077 N38078 10
D38078 N38078 0 diode
R38079 N38078 N38079 10
D38079 N38079 0 diode
R38080 N38079 N38080 10
D38080 N38080 0 diode
R38081 N38080 N38081 10
D38081 N38081 0 diode
R38082 N38081 N38082 10
D38082 N38082 0 diode
R38083 N38082 N38083 10
D38083 N38083 0 diode
R38084 N38083 N38084 10
D38084 N38084 0 diode
R38085 N38084 N38085 10
D38085 N38085 0 diode
R38086 N38085 N38086 10
D38086 N38086 0 diode
R38087 N38086 N38087 10
D38087 N38087 0 diode
R38088 N38087 N38088 10
D38088 N38088 0 diode
R38089 N38088 N38089 10
D38089 N38089 0 diode
R38090 N38089 N38090 10
D38090 N38090 0 diode
R38091 N38090 N38091 10
D38091 N38091 0 diode
R38092 N38091 N38092 10
D38092 N38092 0 diode
R38093 N38092 N38093 10
D38093 N38093 0 diode
R38094 N38093 N38094 10
D38094 N38094 0 diode
R38095 N38094 N38095 10
D38095 N38095 0 diode
R38096 N38095 N38096 10
D38096 N38096 0 diode
R38097 N38096 N38097 10
D38097 N38097 0 diode
R38098 N38097 N38098 10
D38098 N38098 0 diode
R38099 N38098 N38099 10
D38099 N38099 0 diode
R38100 N38099 N38100 10
D38100 N38100 0 diode
R38101 N38100 N38101 10
D38101 N38101 0 diode
R38102 N38101 N38102 10
D38102 N38102 0 diode
R38103 N38102 N38103 10
D38103 N38103 0 diode
R38104 N38103 N38104 10
D38104 N38104 0 diode
R38105 N38104 N38105 10
D38105 N38105 0 diode
R38106 N38105 N38106 10
D38106 N38106 0 diode
R38107 N38106 N38107 10
D38107 N38107 0 diode
R38108 N38107 N38108 10
D38108 N38108 0 diode
R38109 N38108 N38109 10
D38109 N38109 0 diode
R38110 N38109 N38110 10
D38110 N38110 0 diode
R38111 N38110 N38111 10
D38111 N38111 0 diode
R38112 N38111 N38112 10
D38112 N38112 0 diode
R38113 N38112 N38113 10
D38113 N38113 0 diode
R38114 N38113 N38114 10
D38114 N38114 0 diode
R38115 N38114 N38115 10
D38115 N38115 0 diode
R38116 N38115 N38116 10
D38116 N38116 0 diode
R38117 N38116 N38117 10
D38117 N38117 0 diode
R38118 N38117 N38118 10
D38118 N38118 0 diode
R38119 N38118 N38119 10
D38119 N38119 0 diode
R38120 N38119 N38120 10
D38120 N38120 0 diode
R38121 N38120 N38121 10
D38121 N38121 0 diode
R38122 N38121 N38122 10
D38122 N38122 0 diode
R38123 N38122 N38123 10
D38123 N38123 0 diode
R38124 N38123 N38124 10
D38124 N38124 0 diode
R38125 N38124 N38125 10
D38125 N38125 0 diode
R38126 N38125 N38126 10
D38126 N38126 0 diode
R38127 N38126 N38127 10
D38127 N38127 0 diode
R38128 N38127 N38128 10
D38128 N38128 0 diode
R38129 N38128 N38129 10
D38129 N38129 0 diode
R38130 N38129 N38130 10
D38130 N38130 0 diode
R38131 N38130 N38131 10
D38131 N38131 0 diode
R38132 N38131 N38132 10
D38132 N38132 0 diode
R38133 N38132 N38133 10
D38133 N38133 0 diode
R38134 N38133 N38134 10
D38134 N38134 0 diode
R38135 N38134 N38135 10
D38135 N38135 0 diode
R38136 N38135 N38136 10
D38136 N38136 0 diode
R38137 N38136 N38137 10
D38137 N38137 0 diode
R38138 N38137 N38138 10
D38138 N38138 0 diode
R38139 N38138 N38139 10
D38139 N38139 0 diode
R38140 N38139 N38140 10
D38140 N38140 0 diode
R38141 N38140 N38141 10
D38141 N38141 0 diode
R38142 N38141 N38142 10
D38142 N38142 0 diode
R38143 N38142 N38143 10
D38143 N38143 0 diode
R38144 N38143 N38144 10
D38144 N38144 0 diode
R38145 N38144 N38145 10
D38145 N38145 0 diode
R38146 N38145 N38146 10
D38146 N38146 0 diode
R38147 N38146 N38147 10
D38147 N38147 0 diode
R38148 N38147 N38148 10
D38148 N38148 0 diode
R38149 N38148 N38149 10
D38149 N38149 0 diode
R38150 N38149 N38150 10
D38150 N38150 0 diode
R38151 N38150 N38151 10
D38151 N38151 0 diode
R38152 N38151 N38152 10
D38152 N38152 0 diode
R38153 N38152 N38153 10
D38153 N38153 0 diode
R38154 N38153 N38154 10
D38154 N38154 0 diode
R38155 N38154 N38155 10
D38155 N38155 0 diode
R38156 N38155 N38156 10
D38156 N38156 0 diode
R38157 N38156 N38157 10
D38157 N38157 0 diode
R38158 N38157 N38158 10
D38158 N38158 0 diode
R38159 N38158 N38159 10
D38159 N38159 0 diode
R38160 N38159 N38160 10
D38160 N38160 0 diode
R38161 N38160 N38161 10
D38161 N38161 0 diode
R38162 N38161 N38162 10
D38162 N38162 0 diode
R38163 N38162 N38163 10
D38163 N38163 0 diode
R38164 N38163 N38164 10
D38164 N38164 0 diode
R38165 N38164 N38165 10
D38165 N38165 0 diode
R38166 N38165 N38166 10
D38166 N38166 0 diode
R38167 N38166 N38167 10
D38167 N38167 0 diode
R38168 N38167 N38168 10
D38168 N38168 0 diode
R38169 N38168 N38169 10
D38169 N38169 0 diode
R38170 N38169 N38170 10
D38170 N38170 0 diode
R38171 N38170 N38171 10
D38171 N38171 0 diode
R38172 N38171 N38172 10
D38172 N38172 0 diode
R38173 N38172 N38173 10
D38173 N38173 0 diode
R38174 N38173 N38174 10
D38174 N38174 0 diode
R38175 N38174 N38175 10
D38175 N38175 0 diode
R38176 N38175 N38176 10
D38176 N38176 0 diode
R38177 N38176 N38177 10
D38177 N38177 0 diode
R38178 N38177 N38178 10
D38178 N38178 0 diode
R38179 N38178 N38179 10
D38179 N38179 0 diode
R38180 N38179 N38180 10
D38180 N38180 0 diode
R38181 N38180 N38181 10
D38181 N38181 0 diode
R38182 N38181 N38182 10
D38182 N38182 0 diode
R38183 N38182 N38183 10
D38183 N38183 0 diode
R38184 N38183 N38184 10
D38184 N38184 0 diode
R38185 N38184 N38185 10
D38185 N38185 0 diode
R38186 N38185 N38186 10
D38186 N38186 0 diode
R38187 N38186 N38187 10
D38187 N38187 0 diode
R38188 N38187 N38188 10
D38188 N38188 0 diode
R38189 N38188 N38189 10
D38189 N38189 0 diode
R38190 N38189 N38190 10
D38190 N38190 0 diode
R38191 N38190 N38191 10
D38191 N38191 0 diode
R38192 N38191 N38192 10
D38192 N38192 0 diode
R38193 N38192 N38193 10
D38193 N38193 0 diode
R38194 N38193 N38194 10
D38194 N38194 0 diode
R38195 N38194 N38195 10
D38195 N38195 0 diode
R38196 N38195 N38196 10
D38196 N38196 0 diode
R38197 N38196 N38197 10
D38197 N38197 0 diode
R38198 N38197 N38198 10
D38198 N38198 0 diode
R38199 N38198 N38199 10
D38199 N38199 0 diode
R38200 N38199 N38200 10
D38200 N38200 0 diode
R38201 N38200 N38201 10
D38201 N38201 0 diode
R38202 N38201 N38202 10
D38202 N38202 0 diode
R38203 N38202 N38203 10
D38203 N38203 0 diode
R38204 N38203 N38204 10
D38204 N38204 0 diode
R38205 N38204 N38205 10
D38205 N38205 0 diode
R38206 N38205 N38206 10
D38206 N38206 0 diode
R38207 N38206 N38207 10
D38207 N38207 0 diode
R38208 N38207 N38208 10
D38208 N38208 0 diode
R38209 N38208 N38209 10
D38209 N38209 0 diode
R38210 N38209 N38210 10
D38210 N38210 0 diode
R38211 N38210 N38211 10
D38211 N38211 0 diode
R38212 N38211 N38212 10
D38212 N38212 0 diode
R38213 N38212 N38213 10
D38213 N38213 0 diode
R38214 N38213 N38214 10
D38214 N38214 0 diode
R38215 N38214 N38215 10
D38215 N38215 0 diode
R38216 N38215 N38216 10
D38216 N38216 0 diode
R38217 N38216 N38217 10
D38217 N38217 0 diode
R38218 N38217 N38218 10
D38218 N38218 0 diode
R38219 N38218 N38219 10
D38219 N38219 0 diode
R38220 N38219 N38220 10
D38220 N38220 0 diode
R38221 N38220 N38221 10
D38221 N38221 0 diode
R38222 N38221 N38222 10
D38222 N38222 0 diode
R38223 N38222 N38223 10
D38223 N38223 0 diode
R38224 N38223 N38224 10
D38224 N38224 0 diode
R38225 N38224 N38225 10
D38225 N38225 0 diode
R38226 N38225 N38226 10
D38226 N38226 0 diode
R38227 N38226 N38227 10
D38227 N38227 0 diode
R38228 N38227 N38228 10
D38228 N38228 0 diode
R38229 N38228 N38229 10
D38229 N38229 0 diode
R38230 N38229 N38230 10
D38230 N38230 0 diode
R38231 N38230 N38231 10
D38231 N38231 0 diode
R38232 N38231 N38232 10
D38232 N38232 0 diode
R38233 N38232 N38233 10
D38233 N38233 0 diode
R38234 N38233 N38234 10
D38234 N38234 0 diode
R38235 N38234 N38235 10
D38235 N38235 0 diode
R38236 N38235 N38236 10
D38236 N38236 0 diode
R38237 N38236 N38237 10
D38237 N38237 0 diode
R38238 N38237 N38238 10
D38238 N38238 0 diode
R38239 N38238 N38239 10
D38239 N38239 0 diode
R38240 N38239 N38240 10
D38240 N38240 0 diode
R38241 N38240 N38241 10
D38241 N38241 0 diode
R38242 N38241 N38242 10
D38242 N38242 0 diode
R38243 N38242 N38243 10
D38243 N38243 0 diode
R38244 N38243 N38244 10
D38244 N38244 0 diode
R38245 N38244 N38245 10
D38245 N38245 0 diode
R38246 N38245 N38246 10
D38246 N38246 0 diode
R38247 N38246 N38247 10
D38247 N38247 0 diode
R38248 N38247 N38248 10
D38248 N38248 0 diode
R38249 N38248 N38249 10
D38249 N38249 0 diode
R38250 N38249 N38250 10
D38250 N38250 0 diode
R38251 N38250 N38251 10
D38251 N38251 0 diode
R38252 N38251 N38252 10
D38252 N38252 0 diode
R38253 N38252 N38253 10
D38253 N38253 0 diode
R38254 N38253 N38254 10
D38254 N38254 0 diode
R38255 N38254 N38255 10
D38255 N38255 0 diode
R38256 N38255 N38256 10
D38256 N38256 0 diode
R38257 N38256 N38257 10
D38257 N38257 0 diode
R38258 N38257 N38258 10
D38258 N38258 0 diode
R38259 N38258 N38259 10
D38259 N38259 0 diode
R38260 N38259 N38260 10
D38260 N38260 0 diode
R38261 N38260 N38261 10
D38261 N38261 0 diode
R38262 N38261 N38262 10
D38262 N38262 0 diode
R38263 N38262 N38263 10
D38263 N38263 0 diode
R38264 N38263 N38264 10
D38264 N38264 0 diode
R38265 N38264 N38265 10
D38265 N38265 0 diode
R38266 N38265 N38266 10
D38266 N38266 0 diode
R38267 N38266 N38267 10
D38267 N38267 0 diode
R38268 N38267 N38268 10
D38268 N38268 0 diode
R38269 N38268 N38269 10
D38269 N38269 0 diode
R38270 N38269 N38270 10
D38270 N38270 0 diode
R38271 N38270 N38271 10
D38271 N38271 0 diode
R38272 N38271 N38272 10
D38272 N38272 0 diode
R38273 N38272 N38273 10
D38273 N38273 0 diode
R38274 N38273 N38274 10
D38274 N38274 0 diode
R38275 N38274 N38275 10
D38275 N38275 0 diode
R38276 N38275 N38276 10
D38276 N38276 0 diode
R38277 N38276 N38277 10
D38277 N38277 0 diode
R38278 N38277 N38278 10
D38278 N38278 0 diode
R38279 N38278 N38279 10
D38279 N38279 0 diode
R38280 N38279 N38280 10
D38280 N38280 0 diode
R38281 N38280 N38281 10
D38281 N38281 0 diode
R38282 N38281 N38282 10
D38282 N38282 0 diode
R38283 N38282 N38283 10
D38283 N38283 0 diode
R38284 N38283 N38284 10
D38284 N38284 0 diode
R38285 N38284 N38285 10
D38285 N38285 0 diode
R38286 N38285 N38286 10
D38286 N38286 0 diode
R38287 N38286 N38287 10
D38287 N38287 0 diode
R38288 N38287 N38288 10
D38288 N38288 0 diode
R38289 N38288 N38289 10
D38289 N38289 0 diode
R38290 N38289 N38290 10
D38290 N38290 0 diode
R38291 N38290 N38291 10
D38291 N38291 0 diode
R38292 N38291 N38292 10
D38292 N38292 0 diode
R38293 N38292 N38293 10
D38293 N38293 0 diode
R38294 N38293 N38294 10
D38294 N38294 0 diode
R38295 N38294 N38295 10
D38295 N38295 0 diode
R38296 N38295 N38296 10
D38296 N38296 0 diode
R38297 N38296 N38297 10
D38297 N38297 0 diode
R38298 N38297 N38298 10
D38298 N38298 0 diode
R38299 N38298 N38299 10
D38299 N38299 0 diode
R38300 N38299 N38300 10
D38300 N38300 0 diode
R38301 N38300 N38301 10
D38301 N38301 0 diode
R38302 N38301 N38302 10
D38302 N38302 0 diode
R38303 N38302 N38303 10
D38303 N38303 0 diode
R38304 N38303 N38304 10
D38304 N38304 0 diode
R38305 N38304 N38305 10
D38305 N38305 0 diode
R38306 N38305 N38306 10
D38306 N38306 0 diode
R38307 N38306 N38307 10
D38307 N38307 0 diode
R38308 N38307 N38308 10
D38308 N38308 0 diode
R38309 N38308 N38309 10
D38309 N38309 0 diode
R38310 N38309 N38310 10
D38310 N38310 0 diode
R38311 N38310 N38311 10
D38311 N38311 0 diode
R38312 N38311 N38312 10
D38312 N38312 0 diode
R38313 N38312 N38313 10
D38313 N38313 0 diode
R38314 N38313 N38314 10
D38314 N38314 0 diode
R38315 N38314 N38315 10
D38315 N38315 0 diode
R38316 N38315 N38316 10
D38316 N38316 0 diode
R38317 N38316 N38317 10
D38317 N38317 0 diode
R38318 N38317 N38318 10
D38318 N38318 0 diode
R38319 N38318 N38319 10
D38319 N38319 0 diode
R38320 N38319 N38320 10
D38320 N38320 0 diode
R38321 N38320 N38321 10
D38321 N38321 0 diode
R38322 N38321 N38322 10
D38322 N38322 0 diode
R38323 N38322 N38323 10
D38323 N38323 0 diode
R38324 N38323 N38324 10
D38324 N38324 0 diode
R38325 N38324 N38325 10
D38325 N38325 0 diode
R38326 N38325 N38326 10
D38326 N38326 0 diode
R38327 N38326 N38327 10
D38327 N38327 0 diode
R38328 N38327 N38328 10
D38328 N38328 0 diode
R38329 N38328 N38329 10
D38329 N38329 0 diode
R38330 N38329 N38330 10
D38330 N38330 0 diode
R38331 N38330 N38331 10
D38331 N38331 0 diode
R38332 N38331 N38332 10
D38332 N38332 0 diode
R38333 N38332 N38333 10
D38333 N38333 0 diode
R38334 N38333 N38334 10
D38334 N38334 0 diode
R38335 N38334 N38335 10
D38335 N38335 0 diode
R38336 N38335 N38336 10
D38336 N38336 0 diode
R38337 N38336 N38337 10
D38337 N38337 0 diode
R38338 N38337 N38338 10
D38338 N38338 0 diode
R38339 N38338 N38339 10
D38339 N38339 0 diode
R38340 N38339 N38340 10
D38340 N38340 0 diode
R38341 N38340 N38341 10
D38341 N38341 0 diode
R38342 N38341 N38342 10
D38342 N38342 0 diode
R38343 N38342 N38343 10
D38343 N38343 0 diode
R38344 N38343 N38344 10
D38344 N38344 0 diode
R38345 N38344 N38345 10
D38345 N38345 0 diode
R38346 N38345 N38346 10
D38346 N38346 0 diode
R38347 N38346 N38347 10
D38347 N38347 0 diode
R38348 N38347 N38348 10
D38348 N38348 0 diode
R38349 N38348 N38349 10
D38349 N38349 0 diode
R38350 N38349 N38350 10
D38350 N38350 0 diode
R38351 N38350 N38351 10
D38351 N38351 0 diode
R38352 N38351 N38352 10
D38352 N38352 0 diode
R38353 N38352 N38353 10
D38353 N38353 0 diode
R38354 N38353 N38354 10
D38354 N38354 0 diode
R38355 N38354 N38355 10
D38355 N38355 0 diode
R38356 N38355 N38356 10
D38356 N38356 0 diode
R38357 N38356 N38357 10
D38357 N38357 0 diode
R38358 N38357 N38358 10
D38358 N38358 0 diode
R38359 N38358 N38359 10
D38359 N38359 0 diode
R38360 N38359 N38360 10
D38360 N38360 0 diode
R38361 N38360 N38361 10
D38361 N38361 0 diode
R38362 N38361 N38362 10
D38362 N38362 0 diode
R38363 N38362 N38363 10
D38363 N38363 0 diode
R38364 N38363 N38364 10
D38364 N38364 0 diode
R38365 N38364 N38365 10
D38365 N38365 0 diode
R38366 N38365 N38366 10
D38366 N38366 0 diode
R38367 N38366 N38367 10
D38367 N38367 0 diode
R38368 N38367 N38368 10
D38368 N38368 0 diode
R38369 N38368 N38369 10
D38369 N38369 0 diode
R38370 N38369 N38370 10
D38370 N38370 0 diode
R38371 N38370 N38371 10
D38371 N38371 0 diode
R38372 N38371 N38372 10
D38372 N38372 0 diode
R38373 N38372 N38373 10
D38373 N38373 0 diode
R38374 N38373 N38374 10
D38374 N38374 0 diode
R38375 N38374 N38375 10
D38375 N38375 0 diode
R38376 N38375 N38376 10
D38376 N38376 0 diode
R38377 N38376 N38377 10
D38377 N38377 0 diode
R38378 N38377 N38378 10
D38378 N38378 0 diode
R38379 N38378 N38379 10
D38379 N38379 0 diode
R38380 N38379 N38380 10
D38380 N38380 0 diode
R38381 N38380 N38381 10
D38381 N38381 0 diode
R38382 N38381 N38382 10
D38382 N38382 0 diode
R38383 N38382 N38383 10
D38383 N38383 0 diode
R38384 N38383 N38384 10
D38384 N38384 0 diode
R38385 N38384 N38385 10
D38385 N38385 0 diode
R38386 N38385 N38386 10
D38386 N38386 0 diode
R38387 N38386 N38387 10
D38387 N38387 0 diode
R38388 N38387 N38388 10
D38388 N38388 0 diode
R38389 N38388 N38389 10
D38389 N38389 0 diode
R38390 N38389 N38390 10
D38390 N38390 0 diode
R38391 N38390 N38391 10
D38391 N38391 0 diode
R38392 N38391 N38392 10
D38392 N38392 0 diode
R38393 N38392 N38393 10
D38393 N38393 0 diode
R38394 N38393 N38394 10
D38394 N38394 0 diode
R38395 N38394 N38395 10
D38395 N38395 0 diode
R38396 N38395 N38396 10
D38396 N38396 0 diode
R38397 N38396 N38397 10
D38397 N38397 0 diode
R38398 N38397 N38398 10
D38398 N38398 0 diode
R38399 N38398 N38399 10
D38399 N38399 0 diode
R38400 N38399 N38400 10
D38400 N38400 0 diode
R38401 N38400 N38401 10
D38401 N38401 0 diode
R38402 N38401 N38402 10
D38402 N38402 0 diode
R38403 N38402 N38403 10
D38403 N38403 0 diode
R38404 N38403 N38404 10
D38404 N38404 0 diode
R38405 N38404 N38405 10
D38405 N38405 0 diode
R38406 N38405 N38406 10
D38406 N38406 0 diode
R38407 N38406 N38407 10
D38407 N38407 0 diode
R38408 N38407 N38408 10
D38408 N38408 0 diode
R38409 N38408 N38409 10
D38409 N38409 0 diode
R38410 N38409 N38410 10
D38410 N38410 0 diode
R38411 N38410 N38411 10
D38411 N38411 0 diode
R38412 N38411 N38412 10
D38412 N38412 0 diode
R38413 N38412 N38413 10
D38413 N38413 0 diode
R38414 N38413 N38414 10
D38414 N38414 0 diode
R38415 N38414 N38415 10
D38415 N38415 0 diode
R38416 N38415 N38416 10
D38416 N38416 0 diode
R38417 N38416 N38417 10
D38417 N38417 0 diode
R38418 N38417 N38418 10
D38418 N38418 0 diode
R38419 N38418 N38419 10
D38419 N38419 0 diode
R38420 N38419 N38420 10
D38420 N38420 0 diode
R38421 N38420 N38421 10
D38421 N38421 0 diode
R38422 N38421 N38422 10
D38422 N38422 0 diode
R38423 N38422 N38423 10
D38423 N38423 0 diode
R38424 N38423 N38424 10
D38424 N38424 0 diode
R38425 N38424 N38425 10
D38425 N38425 0 diode
R38426 N38425 N38426 10
D38426 N38426 0 diode
R38427 N38426 N38427 10
D38427 N38427 0 diode
R38428 N38427 N38428 10
D38428 N38428 0 diode
R38429 N38428 N38429 10
D38429 N38429 0 diode
R38430 N38429 N38430 10
D38430 N38430 0 diode
R38431 N38430 N38431 10
D38431 N38431 0 diode
R38432 N38431 N38432 10
D38432 N38432 0 diode
R38433 N38432 N38433 10
D38433 N38433 0 diode
R38434 N38433 N38434 10
D38434 N38434 0 diode
R38435 N38434 N38435 10
D38435 N38435 0 diode
R38436 N38435 N38436 10
D38436 N38436 0 diode
R38437 N38436 N38437 10
D38437 N38437 0 diode
R38438 N38437 N38438 10
D38438 N38438 0 diode
R38439 N38438 N38439 10
D38439 N38439 0 diode
R38440 N38439 N38440 10
D38440 N38440 0 diode
R38441 N38440 N38441 10
D38441 N38441 0 diode
R38442 N38441 N38442 10
D38442 N38442 0 diode
R38443 N38442 N38443 10
D38443 N38443 0 diode
R38444 N38443 N38444 10
D38444 N38444 0 diode
R38445 N38444 N38445 10
D38445 N38445 0 diode
R38446 N38445 N38446 10
D38446 N38446 0 diode
R38447 N38446 N38447 10
D38447 N38447 0 diode
R38448 N38447 N38448 10
D38448 N38448 0 diode
R38449 N38448 N38449 10
D38449 N38449 0 diode
R38450 N38449 N38450 10
D38450 N38450 0 diode
R38451 N38450 N38451 10
D38451 N38451 0 diode
R38452 N38451 N38452 10
D38452 N38452 0 diode
R38453 N38452 N38453 10
D38453 N38453 0 diode
R38454 N38453 N38454 10
D38454 N38454 0 diode
R38455 N38454 N38455 10
D38455 N38455 0 diode
R38456 N38455 N38456 10
D38456 N38456 0 diode
R38457 N38456 N38457 10
D38457 N38457 0 diode
R38458 N38457 N38458 10
D38458 N38458 0 diode
R38459 N38458 N38459 10
D38459 N38459 0 diode
R38460 N38459 N38460 10
D38460 N38460 0 diode
R38461 N38460 N38461 10
D38461 N38461 0 diode
R38462 N38461 N38462 10
D38462 N38462 0 diode
R38463 N38462 N38463 10
D38463 N38463 0 diode
R38464 N38463 N38464 10
D38464 N38464 0 diode
R38465 N38464 N38465 10
D38465 N38465 0 diode
R38466 N38465 N38466 10
D38466 N38466 0 diode
R38467 N38466 N38467 10
D38467 N38467 0 diode
R38468 N38467 N38468 10
D38468 N38468 0 diode
R38469 N38468 N38469 10
D38469 N38469 0 diode
R38470 N38469 N38470 10
D38470 N38470 0 diode
R38471 N38470 N38471 10
D38471 N38471 0 diode
R38472 N38471 N38472 10
D38472 N38472 0 diode
R38473 N38472 N38473 10
D38473 N38473 0 diode
R38474 N38473 N38474 10
D38474 N38474 0 diode
R38475 N38474 N38475 10
D38475 N38475 0 diode
R38476 N38475 N38476 10
D38476 N38476 0 diode
R38477 N38476 N38477 10
D38477 N38477 0 diode
R38478 N38477 N38478 10
D38478 N38478 0 diode
R38479 N38478 N38479 10
D38479 N38479 0 diode
R38480 N38479 N38480 10
D38480 N38480 0 diode
R38481 N38480 N38481 10
D38481 N38481 0 diode
R38482 N38481 N38482 10
D38482 N38482 0 diode
R38483 N38482 N38483 10
D38483 N38483 0 diode
R38484 N38483 N38484 10
D38484 N38484 0 diode
R38485 N38484 N38485 10
D38485 N38485 0 diode
R38486 N38485 N38486 10
D38486 N38486 0 diode
R38487 N38486 N38487 10
D38487 N38487 0 diode
R38488 N38487 N38488 10
D38488 N38488 0 diode
R38489 N38488 N38489 10
D38489 N38489 0 diode
R38490 N38489 N38490 10
D38490 N38490 0 diode
R38491 N38490 N38491 10
D38491 N38491 0 diode
R38492 N38491 N38492 10
D38492 N38492 0 diode
R38493 N38492 N38493 10
D38493 N38493 0 diode
R38494 N38493 N38494 10
D38494 N38494 0 diode
R38495 N38494 N38495 10
D38495 N38495 0 diode
R38496 N38495 N38496 10
D38496 N38496 0 diode
R38497 N38496 N38497 10
D38497 N38497 0 diode
R38498 N38497 N38498 10
D38498 N38498 0 diode
R38499 N38498 N38499 10
D38499 N38499 0 diode
R38500 N38499 N38500 10
D38500 N38500 0 diode
R38501 N38500 N38501 10
D38501 N38501 0 diode
R38502 N38501 N38502 10
D38502 N38502 0 diode
R38503 N38502 N38503 10
D38503 N38503 0 diode
R38504 N38503 N38504 10
D38504 N38504 0 diode
R38505 N38504 N38505 10
D38505 N38505 0 diode
R38506 N38505 N38506 10
D38506 N38506 0 diode
R38507 N38506 N38507 10
D38507 N38507 0 diode
R38508 N38507 N38508 10
D38508 N38508 0 diode
R38509 N38508 N38509 10
D38509 N38509 0 diode
R38510 N38509 N38510 10
D38510 N38510 0 diode
R38511 N38510 N38511 10
D38511 N38511 0 diode
R38512 N38511 N38512 10
D38512 N38512 0 diode
R38513 N38512 N38513 10
D38513 N38513 0 diode
R38514 N38513 N38514 10
D38514 N38514 0 diode
R38515 N38514 N38515 10
D38515 N38515 0 diode
R38516 N38515 N38516 10
D38516 N38516 0 diode
R38517 N38516 N38517 10
D38517 N38517 0 diode
R38518 N38517 N38518 10
D38518 N38518 0 diode
R38519 N38518 N38519 10
D38519 N38519 0 diode
R38520 N38519 N38520 10
D38520 N38520 0 diode
R38521 N38520 N38521 10
D38521 N38521 0 diode
R38522 N38521 N38522 10
D38522 N38522 0 diode
R38523 N38522 N38523 10
D38523 N38523 0 diode
R38524 N38523 N38524 10
D38524 N38524 0 diode
R38525 N38524 N38525 10
D38525 N38525 0 diode
R38526 N38525 N38526 10
D38526 N38526 0 diode
R38527 N38526 N38527 10
D38527 N38527 0 diode
R38528 N38527 N38528 10
D38528 N38528 0 diode
R38529 N38528 N38529 10
D38529 N38529 0 diode
R38530 N38529 N38530 10
D38530 N38530 0 diode
R38531 N38530 N38531 10
D38531 N38531 0 diode
R38532 N38531 N38532 10
D38532 N38532 0 diode
R38533 N38532 N38533 10
D38533 N38533 0 diode
R38534 N38533 N38534 10
D38534 N38534 0 diode
R38535 N38534 N38535 10
D38535 N38535 0 diode
R38536 N38535 N38536 10
D38536 N38536 0 diode
R38537 N38536 N38537 10
D38537 N38537 0 diode
R38538 N38537 N38538 10
D38538 N38538 0 diode
R38539 N38538 N38539 10
D38539 N38539 0 diode
R38540 N38539 N38540 10
D38540 N38540 0 diode
R38541 N38540 N38541 10
D38541 N38541 0 diode
R38542 N38541 N38542 10
D38542 N38542 0 diode
R38543 N38542 N38543 10
D38543 N38543 0 diode
R38544 N38543 N38544 10
D38544 N38544 0 diode
R38545 N38544 N38545 10
D38545 N38545 0 diode
R38546 N38545 N38546 10
D38546 N38546 0 diode
R38547 N38546 N38547 10
D38547 N38547 0 diode
R38548 N38547 N38548 10
D38548 N38548 0 diode
R38549 N38548 N38549 10
D38549 N38549 0 diode
R38550 N38549 N38550 10
D38550 N38550 0 diode
R38551 N38550 N38551 10
D38551 N38551 0 diode
R38552 N38551 N38552 10
D38552 N38552 0 diode
R38553 N38552 N38553 10
D38553 N38553 0 diode
R38554 N38553 N38554 10
D38554 N38554 0 diode
R38555 N38554 N38555 10
D38555 N38555 0 diode
R38556 N38555 N38556 10
D38556 N38556 0 diode
R38557 N38556 N38557 10
D38557 N38557 0 diode
R38558 N38557 N38558 10
D38558 N38558 0 diode
R38559 N38558 N38559 10
D38559 N38559 0 diode
R38560 N38559 N38560 10
D38560 N38560 0 diode
R38561 N38560 N38561 10
D38561 N38561 0 diode
R38562 N38561 N38562 10
D38562 N38562 0 diode
R38563 N38562 N38563 10
D38563 N38563 0 diode
R38564 N38563 N38564 10
D38564 N38564 0 diode
R38565 N38564 N38565 10
D38565 N38565 0 diode
R38566 N38565 N38566 10
D38566 N38566 0 diode
R38567 N38566 N38567 10
D38567 N38567 0 diode
R38568 N38567 N38568 10
D38568 N38568 0 diode
R38569 N38568 N38569 10
D38569 N38569 0 diode
R38570 N38569 N38570 10
D38570 N38570 0 diode
R38571 N38570 N38571 10
D38571 N38571 0 diode
R38572 N38571 N38572 10
D38572 N38572 0 diode
R38573 N38572 N38573 10
D38573 N38573 0 diode
R38574 N38573 N38574 10
D38574 N38574 0 diode
R38575 N38574 N38575 10
D38575 N38575 0 diode
R38576 N38575 N38576 10
D38576 N38576 0 diode
R38577 N38576 N38577 10
D38577 N38577 0 diode
R38578 N38577 N38578 10
D38578 N38578 0 diode
R38579 N38578 N38579 10
D38579 N38579 0 diode
R38580 N38579 N38580 10
D38580 N38580 0 diode
R38581 N38580 N38581 10
D38581 N38581 0 diode
R38582 N38581 N38582 10
D38582 N38582 0 diode
R38583 N38582 N38583 10
D38583 N38583 0 diode
R38584 N38583 N38584 10
D38584 N38584 0 diode
R38585 N38584 N38585 10
D38585 N38585 0 diode
R38586 N38585 N38586 10
D38586 N38586 0 diode
R38587 N38586 N38587 10
D38587 N38587 0 diode
R38588 N38587 N38588 10
D38588 N38588 0 diode
R38589 N38588 N38589 10
D38589 N38589 0 diode
R38590 N38589 N38590 10
D38590 N38590 0 diode
R38591 N38590 N38591 10
D38591 N38591 0 diode
R38592 N38591 N38592 10
D38592 N38592 0 diode
R38593 N38592 N38593 10
D38593 N38593 0 diode
R38594 N38593 N38594 10
D38594 N38594 0 diode
R38595 N38594 N38595 10
D38595 N38595 0 diode
R38596 N38595 N38596 10
D38596 N38596 0 diode
R38597 N38596 N38597 10
D38597 N38597 0 diode
R38598 N38597 N38598 10
D38598 N38598 0 diode
R38599 N38598 N38599 10
D38599 N38599 0 diode
R38600 N38599 N38600 10
D38600 N38600 0 diode
R38601 N38600 N38601 10
D38601 N38601 0 diode
R38602 N38601 N38602 10
D38602 N38602 0 diode
R38603 N38602 N38603 10
D38603 N38603 0 diode
R38604 N38603 N38604 10
D38604 N38604 0 diode
R38605 N38604 N38605 10
D38605 N38605 0 diode
R38606 N38605 N38606 10
D38606 N38606 0 diode
R38607 N38606 N38607 10
D38607 N38607 0 diode
R38608 N38607 N38608 10
D38608 N38608 0 diode
R38609 N38608 N38609 10
D38609 N38609 0 diode
R38610 N38609 N38610 10
D38610 N38610 0 diode
R38611 N38610 N38611 10
D38611 N38611 0 diode
R38612 N38611 N38612 10
D38612 N38612 0 diode
R38613 N38612 N38613 10
D38613 N38613 0 diode
R38614 N38613 N38614 10
D38614 N38614 0 diode
R38615 N38614 N38615 10
D38615 N38615 0 diode
R38616 N38615 N38616 10
D38616 N38616 0 diode
R38617 N38616 N38617 10
D38617 N38617 0 diode
R38618 N38617 N38618 10
D38618 N38618 0 diode
R38619 N38618 N38619 10
D38619 N38619 0 diode
R38620 N38619 N38620 10
D38620 N38620 0 diode
R38621 N38620 N38621 10
D38621 N38621 0 diode
R38622 N38621 N38622 10
D38622 N38622 0 diode
R38623 N38622 N38623 10
D38623 N38623 0 diode
R38624 N38623 N38624 10
D38624 N38624 0 diode
R38625 N38624 N38625 10
D38625 N38625 0 diode
R38626 N38625 N38626 10
D38626 N38626 0 diode
R38627 N38626 N38627 10
D38627 N38627 0 diode
R38628 N38627 N38628 10
D38628 N38628 0 diode
R38629 N38628 N38629 10
D38629 N38629 0 diode
R38630 N38629 N38630 10
D38630 N38630 0 diode
R38631 N38630 N38631 10
D38631 N38631 0 diode
R38632 N38631 N38632 10
D38632 N38632 0 diode
R38633 N38632 N38633 10
D38633 N38633 0 diode
R38634 N38633 N38634 10
D38634 N38634 0 diode
R38635 N38634 N38635 10
D38635 N38635 0 diode
R38636 N38635 N38636 10
D38636 N38636 0 diode
R38637 N38636 N38637 10
D38637 N38637 0 diode
R38638 N38637 N38638 10
D38638 N38638 0 diode
R38639 N38638 N38639 10
D38639 N38639 0 diode
R38640 N38639 N38640 10
D38640 N38640 0 diode
R38641 N38640 N38641 10
D38641 N38641 0 diode
R38642 N38641 N38642 10
D38642 N38642 0 diode
R38643 N38642 N38643 10
D38643 N38643 0 diode
R38644 N38643 N38644 10
D38644 N38644 0 diode
R38645 N38644 N38645 10
D38645 N38645 0 diode
R38646 N38645 N38646 10
D38646 N38646 0 diode
R38647 N38646 N38647 10
D38647 N38647 0 diode
R38648 N38647 N38648 10
D38648 N38648 0 diode
R38649 N38648 N38649 10
D38649 N38649 0 diode
R38650 N38649 N38650 10
D38650 N38650 0 diode
R38651 N38650 N38651 10
D38651 N38651 0 diode
R38652 N38651 N38652 10
D38652 N38652 0 diode
R38653 N38652 N38653 10
D38653 N38653 0 diode
R38654 N38653 N38654 10
D38654 N38654 0 diode
R38655 N38654 N38655 10
D38655 N38655 0 diode
R38656 N38655 N38656 10
D38656 N38656 0 diode
R38657 N38656 N38657 10
D38657 N38657 0 diode
R38658 N38657 N38658 10
D38658 N38658 0 diode
R38659 N38658 N38659 10
D38659 N38659 0 diode
R38660 N38659 N38660 10
D38660 N38660 0 diode
R38661 N38660 N38661 10
D38661 N38661 0 diode
R38662 N38661 N38662 10
D38662 N38662 0 diode
R38663 N38662 N38663 10
D38663 N38663 0 diode
R38664 N38663 N38664 10
D38664 N38664 0 diode
R38665 N38664 N38665 10
D38665 N38665 0 diode
R38666 N38665 N38666 10
D38666 N38666 0 diode
R38667 N38666 N38667 10
D38667 N38667 0 diode
R38668 N38667 N38668 10
D38668 N38668 0 diode
R38669 N38668 N38669 10
D38669 N38669 0 diode
R38670 N38669 N38670 10
D38670 N38670 0 diode
R38671 N38670 N38671 10
D38671 N38671 0 diode
R38672 N38671 N38672 10
D38672 N38672 0 diode
R38673 N38672 N38673 10
D38673 N38673 0 diode
R38674 N38673 N38674 10
D38674 N38674 0 diode
R38675 N38674 N38675 10
D38675 N38675 0 diode
R38676 N38675 N38676 10
D38676 N38676 0 diode
R38677 N38676 N38677 10
D38677 N38677 0 diode
R38678 N38677 N38678 10
D38678 N38678 0 diode
R38679 N38678 N38679 10
D38679 N38679 0 diode
R38680 N38679 N38680 10
D38680 N38680 0 diode
R38681 N38680 N38681 10
D38681 N38681 0 diode
R38682 N38681 N38682 10
D38682 N38682 0 diode
R38683 N38682 N38683 10
D38683 N38683 0 diode
R38684 N38683 N38684 10
D38684 N38684 0 diode
R38685 N38684 N38685 10
D38685 N38685 0 diode
R38686 N38685 N38686 10
D38686 N38686 0 diode
R38687 N38686 N38687 10
D38687 N38687 0 diode
R38688 N38687 N38688 10
D38688 N38688 0 diode
R38689 N38688 N38689 10
D38689 N38689 0 diode
R38690 N38689 N38690 10
D38690 N38690 0 diode
R38691 N38690 N38691 10
D38691 N38691 0 diode
R38692 N38691 N38692 10
D38692 N38692 0 diode
R38693 N38692 N38693 10
D38693 N38693 0 diode
R38694 N38693 N38694 10
D38694 N38694 0 diode
R38695 N38694 N38695 10
D38695 N38695 0 diode
R38696 N38695 N38696 10
D38696 N38696 0 diode
R38697 N38696 N38697 10
D38697 N38697 0 diode
R38698 N38697 N38698 10
D38698 N38698 0 diode
R38699 N38698 N38699 10
D38699 N38699 0 diode
R38700 N38699 N38700 10
D38700 N38700 0 diode
R38701 N38700 N38701 10
D38701 N38701 0 diode
R38702 N38701 N38702 10
D38702 N38702 0 diode
R38703 N38702 N38703 10
D38703 N38703 0 diode
R38704 N38703 N38704 10
D38704 N38704 0 diode
R38705 N38704 N38705 10
D38705 N38705 0 diode
R38706 N38705 N38706 10
D38706 N38706 0 diode
R38707 N38706 N38707 10
D38707 N38707 0 diode
R38708 N38707 N38708 10
D38708 N38708 0 diode
R38709 N38708 N38709 10
D38709 N38709 0 diode
R38710 N38709 N38710 10
D38710 N38710 0 diode
R38711 N38710 N38711 10
D38711 N38711 0 diode
R38712 N38711 N38712 10
D38712 N38712 0 diode
R38713 N38712 N38713 10
D38713 N38713 0 diode
R38714 N38713 N38714 10
D38714 N38714 0 diode
R38715 N38714 N38715 10
D38715 N38715 0 diode
R38716 N38715 N38716 10
D38716 N38716 0 diode
R38717 N38716 N38717 10
D38717 N38717 0 diode
R38718 N38717 N38718 10
D38718 N38718 0 diode
R38719 N38718 N38719 10
D38719 N38719 0 diode
R38720 N38719 N38720 10
D38720 N38720 0 diode
R38721 N38720 N38721 10
D38721 N38721 0 diode
R38722 N38721 N38722 10
D38722 N38722 0 diode
R38723 N38722 N38723 10
D38723 N38723 0 diode
R38724 N38723 N38724 10
D38724 N38724 0 diode
R38725 N38724 N38725 10
D38725 N38725 0 diode
R38726 N38725 N38726 10
D38726 N38726 0 diode
R38727 N38726 N38727 10
D38727 N38727 0 diode
R38728 N38727 N38728 10
D38728 N38728 0 diode
R38729 N38728 N38729 10
D38729 N38729 0 diode
R38730 N38729 N38730 10
D38730 N38730 0 diode
R38731 N38730 N38731 10
D38731 N38731 0 diode
R38732 N38731 N38732 10
D38732 N38732 0 diode
R38733 N38732 N38733 10
D38733 N38733 0 diode
R38734 N38733 N38734 10
D38734 N38734 0 diode
R38735 N38734 N38735 10
D38735 N38735 0 diode
R38736 N38735 N38736 10
D38736 N38736 0 diode
R38737 N38736 N38737 10
D38737 N38737 0 diode
R38738 N38737 N38738 10
D38738 N38738 0 diode
R38739 N38738 N38739 10
D38739 N38739 0 diode
R38740 N38739 N38740 10
D38740 N38740 0 diode
R38741 N38740 N38741 10
D38741 N38741 0 diode
R38742 N38741 N38742 10
D38742 N38742 0 diode
R38743 N38742 N38743 10
D38743 N38743 0 diode
R38744 N38743 N38744 10
D38744 N38744 0 diode
R38745 N38744 N38745 10
D38745 N38745 0 diode
R38746 N38745 N38746 10
D38746 N38746 0 diode
R38747 N38746 N38747 10
D38747 N38747 0 diode
R38748 N38747 N38748 10
D38748 N38748 0 diode
R38749 N38748 N38749 10
D38749 N38749 0 diode
R38750 N38749 N38750 10
D38750 N38750 0 diode
R38751 N38750 N38751 10
D38751 N38751 0 diode
R38752 N38751 N38752 10
D38752 N38752 0 diode
R38753 N38752 N38753 10
D38753 N38753 0 diode
R38754 N38753 N38754 10
D38754 N38754 0 diode
R38755 N38754 N38755 10
D38755 N38755 0 diode
R38756 N38755 N38756 10
D38756 N38756 0 diode
R38757 N38756 N38757 10
D38757 N38757 0 diode
R38758 N38757 N38758 10
D38758 N38758 0 diode
R38759 N38758 N38759 10
D38759 N38759 0 diode
R38760 N38759 N38760 10
D38760 N38760 0 diode
R38761 N38760 N38761 10
D38761 N38761 0 diode
R38762 N38761 N38762 10
D38762 N38762 0 diode
R38763 N38762 N38763 10
D38763 N38763 0 diode
R38764 N38763 N38764 10
D38764 N38764 0 diode
R38765 N38764 N38765 10
D38765 N38765 0 diode
R38766 N38765 N38766 10
D38766 N38766 0 diode
R38767 N38766 N38767 10
D38767 N38767 0 diode
R38768 N38767 N38768 10
D38768 N38768 0 diode
R38769 N38768 N38769 10
D38769 N38769 0 diode
R38770 N38769 N38770 10
D38770 N38770 0 diode
R38771 N38770 N38771 10
D38771 N38771 0 diode
R38772 N38771 N38772 10
D38772 N38772 0 diode
R38773 N38772 N38773 10
D38773 N38773 0 diode
R38774 N38773 N38774 10
D38774 N38774 0 diode
R38775 N38774 N38775 10
D38775 N38775 0 diode
R38776 N38775 N38776 10
D38776 N38776 0 diode
R38777 N38776 N38777 10
D38777 N38777 0 diode
R38778 N38777 N38778 10
D38778 N38778 0 diode
R38779 N38778 N38779 10
D38779 N38779 0 diode
R38780 N38779 N38780 10
D38780 N38780 0 diode
R38781 N38780 N38781 10
D38781 N38781 0 diode
R38782 N38781 N38782 10
D38782 N38782 0 diode
R38783 N38782 N38783 10
D38783 N38783 0 diode
R38784 N38783 N38784 10
D38784 N38784 0 diode
R38785 N38784 N38785 10
D38785 N38785 0 diode
R38786 N38785 N38786 10
D38786 N38786 0 diode
R38787 N38786 N38787 10
D38787 N38787 0 diode
R38788 N38787 N38788 10
D38788 N38788 0 diode
R38789 N38788 N38789 10
D38789 N38789 0 diode
R38790 N38789 N38790 10
D38790 N38790 0 diode
R38791 N38790 N38791 10
D38791 N38791 0 diode
R38792 N38791 N38792 10
D38792 N38792 0 diode
R38793 N38792 N38793 10
D38793 N38793 0 diode
R38794 N38793 N38794 10
D38794 N38794 0 diode
R38795 N38794 N38795 10
D38795 N38795 0 diode
R38796 N38795 N38796 10
D38796 N38796 0 diode
R38797 N38796 N38797 10
D38797 N38797 0 diode
R38798 N38797 N38798 10
D38798 N38798 0 diode
R38799 N38798 N38799 10
D38799 N38799 0 diode
R38800 N38799 N38800 10
D38800 N38800 0 diode
R38801 N38800 N38801 10
D38801 N38801 0 diode
R38802 N38801 N38802 10
D38802 N38802 0 diode
R38803 N38802 N38803 10
D38803 N38803 0 diode
R38804 N38803 N38804 10
D38804 N38804 0 diode
R38805 N38804 N38805 10
D38805 N38805 0 diode
R38806 N38805 N38806 10
D38806 N38806 0 diode
R38807 N38806 N38807 10
D38807 N38807 0 diode
R38808 N38807 N38808 10
D38808 N38808 0 diode
R38809 N38808 N38809 10
D38809 N38809 0 diode
R38810 N38809 N38810 10
D38810 N38810 0 diode
R38811 N38810 N38811 10
D38811 N38811 0 diode
R38812 N38811 N38812 10
D38812 N38812 0 diode
R38813 N38812 N38813 10
D38813 N38813 0 diode
R38814 N38813 N38814 10
D38814 N38814 0 diode
R38815 N38814 N38815 10
D38815 N38815 0 diode
R38816 N38815 N38816 10
D38816 N38816 0 diode
R38817 N38816 N38817 10
D38817 N38817 0 diode
R38818 N38817 N38818 10
D38818 N38818 0 diode
R38819 N38818 N38819 10
D38819 N38819 0 diode
R38820 N38819 N38820 10
D38820 N38820 0 diode
R38821 N38820 N38821 10
D38821 N38821 0 diode
R38822 N38821 N38822 10
D38822 N38822 0 diode
R38823 N38822 N38823 10
D38823 N38823 0 diode
R38824 N38823 N38824 10
D38824 N38824 0 diode
R38825 N38824 N38825 10
D38825 N38825 0 diode
R38826 N38825 N38826 10
D38826 N38826 0 diode
R38827 N38826 N38827 10
D38827 N38827 0 diode
R38828 N38827 N38828 10
D38828 N38828 0 diode
R38829 N38828 N38829 10
D38829 N38829 0 diode
R38830 N38829 N38830 10
D38830 N38830 0 diode
R38831 N38830 N38831 10
D38831 N38831 0 diode
R38832 N38831 N38832 10
D38832 N38832 0 diode
R38833 N38832 N38833 10
D38833 N38833 0 diode
R38834 N38833 N38834 10
D38834 N38834 0 diode
R38835 N38834 N38835 10
D38835 N38835 0 diode
R38836 N38835 N38836 10
D38836 N38836 0 diode
R38837 N38836 N38837 10
D38837 N38837 0 diode
R38838 N38837 N38838 10
D38838 N38838 0 diode
R38839 N38838 N38839 10
D38839 N38839 0 diode
R38840 N38839 N38840 10
D38840 N38840 0 diode
R38841 N38840 N38841 10
D38841 N38841 0 diode
R38842 N38841 N38842 10
D38842 N38842 0 diode
R38843 N38842 N38843 10
D38843 N38843 0 diode
R38844 N38843 N38844 10
D38844 N38844 0 diode
R38845 N38844 N38845 10
D38845 N38845 0 diode
R38846 N38845 N38846 10
D38846 N38846 0 diode
R38847 N38846 N38847 10
D38847 N38847 0 diode
R38848 N38847 N38848 10
D38848 N38848 0 diode
R38849 N38848 N38849 10
D38849 N38849 0 diode
R38850 N38849 N38850 10
D38850 N38850 0 diode
R38851 N38850 N38851 10
D38851 N38851 0 diode
R38852 N38851 N38852 10
D38852 N38852 0 diode
R38853 N38852 N38853 10
D38853 N38853 0 diode
R38854 N38853 N38854 10
D38854 N38854 0 diode
R38855 N38854 N38855 10
D38855 N38855 0 diode
R38856 N38855 N38856 10
D38856 N38856 0 diode
R38857 N38856 N38857 10
D38857 N38857 0 diode
R38858 N38857 N38858 10
D38858 N38858 0 diode
R38859 N38858 N38859 10
D38859 N38859 0 diode
R38860 N38859 N38860 10
D38860 N38860 0 diode
R38861 N38860 N38861 10
D38861 N38861 0 diode
R38862 N38861 N38862 10
D38862 N38862 0 diode
R38863 N38862 N38863 10
D38863 N38863 0 diode
R38864 N38863 N38864 10
D38864 N38864 0 diode
R38865 N38864 N38865 10
D38865 N38865 0 diode
R38866 N38865 N38866 10
D38866 N38866 0 diode
R38867 N38866 N38867 10
D38867 N38867 0 diode
R38868 N38867 N38868 10
D38868 N38868 0 diode
R38869 N38868 N38869 10
D38869 N38869 0 diode
R38870 N38869 N38870 10
D38870 N38870 0 diode
R38871 N38870 N38871 10
D38871 N38871 0 diode
R38872 N38871 N38872 10
D38872 N38872 0 diode
R38873 N38872 N38873 10
D38873 N38873 0 diode
R38874 N38873 N38874 10
D38874 N38874 0 diode
R38875 N38874 N38875 10
D38875 N38875 0 diode
R38876 N38875 N38876 10
D38876 N38876 0 diode
R38877 N38876 N38877 10
D38877 N38877 0 diode
R38878 N38877 N38878 10
D38878 N38878 0 diode
R38879 N38878 N38879 10
D38879 N38879 0 diode
R38880 N38879 N38880 10
D38880 N38880 0 diode
R38881 N38880 N38881 10
D38881 N38881 0 diode
R38882 N38881 N38882 10
D38882 N38882 0 diode
R38883 N38882 N38883 10
D38883 N38883 0 diode
R38884 N38883 N38884 10
D38884 N38884 0 diode
R38885 N38884 N38885 10
D38885 N38885 0 diode
R38886 N38885 N38886 10
D38886 N38886 0 diode
R38887 N38886 N38887 10
D38887 N38887 0 diode
R38888 N38887 N38888 10
D38888 N38888 0 diode
R38889 N38888 N38889 10
D38889 N38889 0 diode
R38890 N38889 N38890 10
D38890 N38890 0 diode
R38891 N38890 N38891 10
D38891 N38891 0 diode
R38892 N38891 N38892 10
D38892 N38892 0 diode
R38893 N38892 N38893 10
D38893 N38893 0 diode
R38894 N38893 N38894 10
D38894 N38894 0 diode
R38895 N38894 N38895 10
D38895 N38895 0 diode
R38896 N38895 N38896 10
D38896 N38896 0 diode
R38897 N38896 N38897 10
D38897 N38897 0 diode
R38898 N38897 N38898 10
D38898 N38898 0 diode
R38899 N38898 N38899 10
D38899 N38899 0 diode
R38900 N38899 N38900 10
D38900 N38900 0 diode
R38901 N38900 N38901 10
D38901 N38901 0 diode
R38902 N38901 N38902 10
D38902 N38902 0 diode
R38903 N38902 N38903 10
D38903 N38903 0 diode
R38904 N38903 N38904 10
D38904 N38904 0 diode
R38905 N38904 N38905 10
D38905 N38905 0 diode
R38906 N38905 N38906 10
D38906 N38906 0 diode
R38907 N38906 N38907 10
D38907 N38907 0 diode
R38908 N38907 N38908 10
D38908 N38908 0 diode
R38909 N38908 N38909 10
D38909 N38909 0 diode
R38910 N38909 N38910 10
D38910 N38910 0 diode
R38911 N38910 N38911 10
D38911 N38911 0 diode
R38912 N38911 N38912 10
D38912 N38912 0 diode
R38913 N38912 N38913 10
D38913 N38913 0 diode
R38914 N38913 N38914 10
D38914 N38914 0 diode
R38915 N38914 N38915 10
D38915 N38915 0 diode
R38916 N38915 N38916 10
D38916 N38916 0 diode
R38917 N38916 N38917 10
D38917 N38917 0 diode
R38918 N38917 N38918 10
D38918 N38918 0 diode
R38919 N38918 N38919 10
D38919 N38919 0 diode
R38920 N38919 N38920 10
D38920 N38920 0 diode
R38921 N38920 N38921 10
D38921 N38921 0 diode
R38922 N38921 N38922 10
D38922 N38922 0 diode
R38923 N38922 N38923 10
D38923 N38923 0 diode
R38924 N38923 N38924 10
D38924 N38924 0 diode
R38925 N38924 N38925 10
D38925 N38925 0 diode
R38926 N38925 N38926 10
D38926 N38926 0 diode
R38927 N38926 N38927 10
D38927 N38927 0 diode
R38928 N38927 N38928 10
D38928 N38928 0 diode
R38929 N38928 N38929 10
D38929 N38929 0 diode
R38930 N38929 N38930 10
D38930 N38930 0 diode
R38931 N38930 N38931 10
D38931 N38931 0 diode
R38932 N38931 N38932 10
D38932 N38932 0 diode
R38933 N38932 N38933 10
D38933 N38933 0 diode
R38934 N38933 N38934 10
D38934 N38934 0 diode
R38935 N38934 N38935 10
D38935 N38935 0 diode
R38936 N38935 N38936 10
D38936 N38936 0 diode
R38937 N38936 N38937 10
D38937 N38937 0 diode
R38938 N38937 N38938 10
D38938 N38938 0 diode
R38939 N38938 N38939 10
D38939 N38939 0 diode
R38940 N38939 N38940 10
D38940 N38940 0 diode
R38941 N38940 N38941 10
D38941 N38941 0 diode
R38942 N38941 N38942 10
D38942 N38942 0 diode
R38943 N38942 N38943 10
D38943 N38943 0 diode
R38944 N38943 N38944 10
D38944 N38944 0 diode
R38945 N38944 N38945 10
D38945 N38945 0 diode
R38946 N38945 N38946 10
D38946 N38946 0 diode
R38947 N38946 N38947 10
D38947 N38947 0 diode
R38948 N38947 N38948 10
D38948 N38948 0 diode
R38949 N38948 N38949 10
D38949 N38949 0 diode
R38950 N38949 N38950 10
D38950 N38950 0 diode
R38951 N38950 N38951 10
D38951 N38951 0 diode
R38952 N38951 N38952 10
D38952 N38952 0 diode
R38953 N38952 N38953 10
D38953 N38953 0 diode
R38954 N38953 N38954 10
D38954 N38954 0 diode
R38955 N38954 N38955 10
D38955 N38955 0 diode
R38956 N38955 N38956 10
D38956 N38956 0 diode
R38957 N38956 N38957 10
D38957 N38957 0 diode
R38958 N38957 N38958 10
D38958 N38958 0 diode
R38959 N38958 N38959 10
D38959 N38959 0 diode
R38960 N38959 N38960 10
D38960 N38960 0 diode
R38961 N38960 N38961 10
D38961 N38961 0 diode
R38962 N38961 N38962 10
D38962 N38962 0 diode
R38963 N38962 N38963 10
D38963 N38963 0 diode
R38964 N38963 N38964 10
D38964 N38964 0 diode
R38965 N38964 N38965 10
D38965 N38965 0 diode
R38966 N38965 N38966 10
D38966 N38966 0 diode
R38967 N38966 N38967 10
D38967 N38967 0 diode
R38968 N38967 N38968 10
D38968 N38968 0 diode
R38969 N38968 N38969 10
D38969 N38969 0 diode
R38970 N38969 N38970 10
D38970 N38970 0 diode
R38971 N38970 N38971 10
D38971 N38971 0 diode
R38972 N38971 N38972 10
D38972 N38972 0 diode
R38973 N38972 N38973 10
D38973 N38973 0 diode
R38974 N38973 N38974 10
D38974 N38974 0 diode
R38975 N38974 N38975 10
D38975 N38975 0 diode
R38976 N38975 N38976 10
D38976 N38976 0 diode
R38977 N38976 N38977 10
D38977 N38977 0 diode
R38978 N38977 N38978 10
D38978 N38978 0 diode
R38979 N38978 N38979 10
D38979 N38979 0 diode
R38980 N38979 N38980 10
D38980 N38980 0 diode
R38981 N38980 N38981 10
D38981 N38981 0 diode
R38982 N38981 N38982 10
D38982 N38982 0 diode
R38983 N38982 N38983 10
D38983 N38983 0 diode
R38984 N38983 N38984 10
D38984 N38984 0 diode
R38985 N38984 N38985 10
D38985 N38985 0 diode
R38986 N38985 N38986 10
D38986 N38986 0 diode
R38987 N38986 N38987 10
D38987 N38987 0 diode
R38988 N38987 N38988 10
D38988 N38988 0 diode
R38989 N38988 N38989 10
D38989 N38989 0 diode
R38990 N38989 N38990 10
D38990 N38990 0 diode
R38991 N38990 N38991 10
D38991 N38991 0 diode
R38992 N38991 N38992 10
D38992 N38992 0 diode
R38993 N38992 N38993 10
D38993 N38993 0 diode
R38994 N38993 N38994 10
D38994 N38994 0 diode
R38995 N38994 N38995 10
D38995 N38995 0 diode
R38996 N38995 N38996 10
D38996 N38996 0 diode
R38997 N38996 N38997 10
D38997 N38997 0 diode
R38998 N38997 N38998 10
D38998 N38998 0 diode
R38999 N38998 N38999 10
D38999 N38999 0 diode
R39000 N38999 N39000 10
D39000 N39000 0 diode
R39001 N39000 N39001 10
D39001 N39001 0 diode
R39002 N39001 N39002 10
D39002 N39002 0 diode
R39003 N39002 N39003 10
D39003 N39003 0 diode
R39004 N39003 N39004 10
D39004 N39004 0 diode
R39005 N39004 N39005 10
D39005 N39005 0 diode
R39006 N39005 N39006 10
D39006 N39006 0 diode
R39007 N39006 N39007 10
D39007 N39007 0 diode
R39008 N39007 N39008 10
D39008 N39008 0 diode
R39009 N39008 N39009 10
D39009 N39009 0 diode
R39010 N39009 N39010 10
D39010 N39010 0 diode
R39011 N39010 N39011 10
D39011 N39011 0 diode
R39012 N39011 N39012 10
D39012 N39012 0 diode
R39013 N39012 N39013 10
D39013 N39013 0 diode
R39014 N39013 N39014 10
D39014 N39014 0 diode
R39015 N39014 N39015 10
D39015 N39015 0 diode
R39016 N39015 N39016 10
D39016 N39016 0 diode
R39017 N39016 N39017 10
D39017 N39017 0 diode
R39018 N39017 N39018 10
D39018 N39018 0 diode
R39019 N39018 N39019 10
D39019 N39019 0 diode
R39020 N39019 N39020 10
D39020 N39020 0 diode
R39021 N39020 N39021 10
D39021 N39021 0 diode
R39022 N39021 N39022 10
D39022 N39022 0 diode
R39023 N39022 N39023 10
D39023 N39023 0 diode
R39024 N39023 N39024 10
D39024 N39024 0 diode
R39025 N39024 N39025 10
D39025 N39025 0 diode
R39026 N39025 N39026 10
D39026 N39026 0 diode
R39027 N39026 N39027 10
D39027 N39027 0 diode
R39028 N39027 N39028 10
D39028 N39028 0 diode
R39029 N39028 N39029 10
D39029 N39029 0 diode
R39030 N39029 N39030 10
D39030 N39030 0 diode
R39031 N39030 N39031 10
D39031 N39031 0 diode
R39032 N39031 N39032 10
D39032 N39032 0 diode
R39033 N39032 N39033 10
D39033 N39033 0 diode
R39034 N39033 N39034 10
D39034 N39034 0 diode
R39035 N39034 N39035 10
D39035 N39035 0 diode
R39036 N39035 N39036 10
D39036 N39036 0 diode
R39037 N39036 N39037 10
D39037 N39037 0 diode
R39038 N39037 N39038 10
D39038 N39038 0 diode
R39039 N39038 N39039 10
D39039 N39039 0 diode
R39040 N39039 N39040 10
D39040 N39040 0 diode
R39041 N39040 N39041 10
D39041 N39041 0 diode
R39042 N39041 N39042 10
D39042 N39042 0 diode
R39043 N39042 N39043 10
D39043 N39043 0 diode
R39044 N39043 N39044 10
D39044 N39044 0 diode
R39045 N39044 N39045 10
D39045 N39045 0 diode
R39046 N39045 N39046 10
D39046 N39046 0 diode
R39047 N39046 N39047 10
D39047 N39047 0 diode
R39048 N39047 N39048 10
D39048 N39048 0 diode
R39049 N39048 N39049 10
D39049 N39049 0 diode
R39050 N39049 N39050 10
D39050 N39050 0 diode
R39051 N39050 N39051 10
D39051 N39051 0 diode
R39052 N39051 N39052 10
D39052 N39052 0 diode
R39053 N39052 N39053 10
D39053 N39053 0 diode
R39054 N39053 N39054 10
D39054 N39054 0 diode
R39055 N39054 N39055 10
D39055 N39055 0 diode
R39056 N39055 N39056 10
D39056 N39056 0 diode
R39057 N39056 N39057 10
D39057 N39057 0 diode
R39058 N39057 N39058 10
D39058 N39058 0 diode
R39059 N39058 N39059 10
D39059 N39059 0 diode
R39060 N39059 N39060 10
D39060 N39060 0 diode
R39061 N39060 N39061 10
D39061 N39061 0 diode
R39062 N39061 N39062 10
D39062 N39062 0 diode
R39063 N39062 N39063 10
D39063 N39063 0 diode
R39064 N39063 N39064 10
D39064 N39064 0 diode
R39065 N39064 N39065 10
D39065 N39065 0 diode
R39066 N39065 N39066 10
D39066 N39066 0 diode
R39067 N39066 N39067 10
D39067 N39067 0 diode
R39068 N39067 N39068 10
D39068 N39068 0 diode
R39069 N39068 N39069 10
D39069 N39069 0 diode
R39070 N39069 N39070 10
D39070 N39070 0 diode
R39071 N39070 N39071 10
D39071 N39071 0 diode
R39072 N39071 N39072 10
D39072 N39072 0 diode
R39073 N39072 N39073 10
D39073 N39073 0 diode
R39074 N39073 N39074 10
D39074 N39074 0 diode
R39075 N39074 N39075 10
D39075 N39075 0 diode
R39076 N39075 N39076 10
D39076 N39076 0 diode
R39077 N39076 N39077 10
D39077 N39077 0 diode
R39078 N39077 N39078 10
D39078 N39078 0 diode
R39079 N39078 N39079 10
D39079 N39079 0 diode
R39080 N39079 N39080 10
D39080 N39080 0 diode
R39081 N39080 N39081 10
D39081 N39081 0 diode
R39082 N39081 N39082 10
D39082 N39082 0 diode
R39083 N39082 N39083 10
D39083 N39083 0 diode
R39084 N39083 N39084 10
D39084 N39084 0 diode
R39085 N39084 N39085 10
D39085 N39085 0 diode
R39086 N39085 N39086 10
D39086 N39086 0 diode
R39087 N39086 N39087 10
D39087 N39087 0 diode
R39088 N39087 N39088 10
D39088 N39088 0 diode
R39089 N39088 N39089 10
D39089 N39089 0 diode
R39090 N39089 N39090 10
D39090 N39090 0 diode
R39091 N39090 N39091 10
D39091 N39091 0 diode
R39092 N39091 N39092 10
D39092 N39092 0 diode
R39093 N39092 N39093 10
D39093 N39093 0 diode
R39094 N39093 N39094 10
D39094 N39094 0 diode
R39095 N39094 N39095 10
D39095 N39095 0 diode
R39096 N39095 N39096 10
D39096 N39096 0 diode
R39097 N39096 N39097 10
D39097 N39097 0 diode
R39098 N39097 N39098 10
D39098 N39098 0 diode
R39099 N39098 N39099 10
D39099 N39099 0 diode
R39100 N39099 N39100 10
D39100 N39100 0 diode
R39101 N39100 N39101 10
D39101 N39101 0 diode
R39102 N39101 N39102 10
D39102 N39102 0 diode
R39103 N39102 N39103 10
D39103 N39103 0 diode
R39104 N39103 N39104 10
D39104 N39104 0 diode
R39105 N39104 N39105 10
D39105 N39105 0 diode
R39106 N39105 N39106 10
D39106 N39106 0 diode
R39107 N39106 N39107 10
D39107 N39107 0 diode
R39108 N39107 N39108 10
D39108 N39108 0 diode
R39109 N39108 N39109 10
D39109 N39109 0 diode
R39110 N39109 N39110 10
D39110 N39110 0 diode
R39111 N39110 N39111 10
D39111 N39111 0 diode
R39112 N39111 N39112 10
D39112 N39112 0 diode
R39113 N39112 N39113 10
D39113 N39113 0 diode
R39114 N39113 N39114 10
D39114 N39114 0 diode
R39115 N39114 N39115 10
D39115 N39115 0 diode
R39116 N39115 N39116 10
D39116 N39116 0 diode
R39117 N39116 N39117 10
D39117 N39117 0 diode
R39118 N39117 N39118 10
D39118 N39118 0 diode
R39119 N39118 N39119 10
D39119 N39119 0 diode
R39120 N39119 N39120 10
D39120 N39120 0 diode
R39121 N39120 N39121 10
D39121 N39121 0 diode
R39122 N39121 N39122 10
D39122 N39122 0 diode
R39123 N39122 N39123 10
D39123 N39123 0 diode
R39124 N39123 N39124 10
D39124 N39124 0 diode
R39125 N39124 N39125 10
D39125 N39125 0 diode
R39126 N39125 N39126 10
D39126 N39126 0 diode
R39127 N39126 N39127 10
D39127 N39127 0 diode
R39128 N39127 N39128 10
D39128 N39128 0 diode
R39129 N39128 N39129 10
D39129 N39129 0 diode
R39130 N39129 N39130 10
D39130 N39130 0 diode
R39131 N39130 N39131 10
D39131 N39131 0 diode
R39132 N39131 N39132 10
D39132 N39132 0 diode
R39133 N39132 N39133 10
D39133 N39133 0 diode
R39134 N39133 N39134 10
D39134 N39134 0 diode
R39135 N39134 N39135 10
D39135 N39135 0 diode
R39136 N39135 N39136 10
D39136 N39136 0 diode
R39137 N39136 N39137 10
D39137 N39137 0 diode
R39138 N39137 N39138 10
D39138 N39138 0 diode
R39139 N39138 N39139 10
D39139 N39139 0 diode
R39140 N39139 N39140 10
D39140 N39140 0 diode
R39141 N39140 N39141 10
D39141 N39141 0 diode
R39142 N39141 N39142 10
D39142 N39142 0 diode
R39143 N39142 N39143 10
D39143 N39143 0 diode
R39144 N39143 N39144 10
D39144 N39144 0 diode
R39145 N39144 N39145 10
D39145 N39145 0 diode
R39146 N39145 N39146 10
D39146 N39146 0 diode
R39147 N39146 N39147 10
D39147 N39147 0 diode
R39148 N39147 N39148 10
D39148 N39148 0 diode
R39149 N39148 N39149 10
D39149 N39149 0 diode
R39150 N39149 N39150 10
D39150 N39150 0 diode
R39151 N39150 N39151 10
D39151 N39151 0 diode
R39152 N39151 N39152 10
D39152 N39152 0 diode
R39153 N39152 N39153 10
D39153 N39153 0 diode
R39154 N39153 N39154 10
D39154 N39154 0 diode
R39155 N39154 N39155 10
D39155 N39155 0 diode
R39156 N39155 N39156 10
D39156 N39156 0 diode
R39157 N39156 N39157 10
D39157 N39157 0 diode
R39158 N39157 N39158 10
D39158 N39158 0 diode
R39159 N39158 N39159 10
D39159 N39159 0 diode
R39160 N39159 N39160 10
D39160 N39160 0 diode
R39161 N39160 N39161 10
D39161 N39161 0 diode
R39162 N39161 N39162 10
D39162 N39162 0 diode
R39163 N39162 N39163 10
D39163 N39163 0 diode
R39164 N39163 N39164 10
D39164 N39164 0 diode
R39165 N39164 N39165 10
D39165 N39165 0 diode
R39166 N39165 N39166 10
D39166 N39166 0 diode
R39167 N39166 N39167 10
D39167 N39167 0 diode
R39168 N39167 N39168 10
D39168 N39168 0 diode
R39169 N39168 N39169 10
D39169 N39169 0 diode
R39170 N39169 N39170 10
D39170 N39170 0 diode
R39171 N39170 N39171 10
D39171 N39171 0 diode
R39172 N39171 N39172 10
D39172 N39172 0 diode
R39173 N39172 N39173 10
D39173 N39173 0 diode
R39174 N39173 N39174 10
D39174 N39174 0 diode
R39175 N39174 N39175 10
D39175 N39175 0 diode
R39176 N39175 N39176 10
D39176 N39176 0 diode
R39177 N39176 N39177 10
D39177 N39177 0 diode
R39178 N39177 N39178 10
D39178 N39178 0 diode
R39179 N39178 N39179 10
D39179 N39179 0 diode
R39180 N39179 N39180 10
D39180 N39180 0 diode
R39181 N39180 N39181 10
D39181 N39181 0 diode
R39182 N39181 N39182 10
D39182 N39182 0 diode
R39183 N39182 N39183 10
D39183 N39183 0 diode
R39184 N39183 N39184 10
D39184 N39184 0 diode
R39185 N39184 N39185 10
D39185 N39185 0 diode
R39186 N39185 N39186 10
D39186 N39186 0 diode
R39187 N39186 N39187 10
D39187 N39187 0 diode
R39188 N39187 N39188 10
D39188 N39188 0 diode
R39189 N39188 N39189 10
D39189 N39189 0 diode
R39190 N39189 N39190 10
D39190 N39190 0 diode
R39191 N39190 N39191 10
D39191 N39191 0 diode
R39192 N39191 N39192 10
D39192 N39192 0 diode
R39193 N39192 N39193 10
D39193 N39193 0 diode
R39194 N39193 N39194 10
D39194 N39194 0 diode
R39195 N39194 N39195 10
D39195 N39195 0 diode
R39196 N39195 N39196 10
D39196 N39196 0 diode
R39197 N39196 N39197 10
D39197 N39197 0 diode
R39198 N39197 N39198 10
D39198 N39198 0 diode
R39199 N39198 N39199 10
D39199 N39199 0 diode
R39200 N39199 N39200 10
D39200 N39200 0 diode
R39201 N39200 N39201 10
D39201 N39201 0 diode
R39202 N39201 N39202 10
D39202 N39202 0 diode
R39203 N39202 N39203 10
D39203 N39203 0 diode
R39204 N39203 N39204 10
D39204 N39204 0 diode
R39205 N39204 N39205 10
D39205 N39205 0 diode
R39206 N39205 N39206 10
D39206 N39206 0 diode
R39207 N39206 N39207 10
D39207 N39207 0 diode
R39208 N39207 N39208 10
D39208 N39208 0 diode
R39209 N39208 N39209 10
D39209 N39209 0 diode
R39210 N39209 N39210 10
D39210 N39210 0 diode
R39211 N39210 N39211 10
D39211 N39211 0 diode
R39212 N39211 N39212 10
D39212 N39212 0 diode
R39213 N39212 N39213 10
D39213 N39213 0 diode
R39214 N39213 N39214 10
D39214 N39214 0 diode
R39215 N39214 N39215 10
D39215 N39215 0 diode
R39216 N39215 N39216 10
D39216 N39216 0 diode
R39217 N39216 N39217 10
D39217 N39217 0 diode
R39218 N39217 N39218 10
D39218 N39218 0 diode
R39219 N39218 N39219 10
D39219 N39219 0 diode
R39220 N39219 N39220 10
D39220 N39220 0 diode
R39221 N39220 N39221 10
D39221 N39221 0 diode
R39222 N39221 N39222 10
D39222 N39222 0 diode
R39223 N39222 N39223 10
D39223 N39223 0 diode
R39224 N39223 N39224 10
D39224 N39224 0 diode
R39225 N39224 N39225 10
D39225 N39225 0 diode
R39226 N39225 N39226 10
D39226 N39226 0 diode
R39227 N39226 N39227 10
D39227 N39227 0 diode
R39228 N39227 N39228 10
D39228 N39228 0 diode
R39229 N39228 N39229 10
D39229 N39229 0 diode
R39230 N39229 N39230 10
D39230 N39230 0 diode
R39231 N39230 N39231 10
D39231 N39231 0 diode
R39232 N39231 N39232 10
D39232 N39232 0 diode
R39233 N39232 N39233 10
D39233 N39233 0 diode
R39234 N39233 N39234 10
D39234 N39234 0 diode
R39235 N39234 N39235 10
D39235 N39235 0 diode
R39236 N39235 N39236 10
D39236 N39236 0 diode
R39237 N39236 N39237 10
D39237 N39237 0 diode
R39238 N39237 N39238 10
D39238 N39238 0 diode
R39239 N39238 N39239 10
D39239 N39239 0 diode
R39240 N39239 N39240 10
D39240 N39240 0 diode
R39241 N39240 N39241 10
D39241 N39241 0 diode
R39242 N39241 N39242 10
D39242 N39242 0 diode
R39243 N39242 N39243 10
D39243 N39243 0 diode
R39244 N39243 N39244 10
D39244 N39244 0 diode
R39245 N39244 N39245 10
D39245 N39245 0 diode
R39246 N39245 N39246 10
D39246 N39246 0 diode
R39247 N39246 N39247 10
D39247 N39247 0 diode
R39248 N39247 N39248 10
D39248 N39248 0 diode
R39249 N39248 N39249 10
D39249 N39249 0 diode
R39250 N39249 N39250 10
D39250 N39250 0 diode
R39251 N39250 N39251 10
D39251 N39251 0 diode
R39252 N39251 N39252 10
D39252 N39252 0 diode
R39253 N39252 N39253 10
D39253 N39253 0 diode
R39254 N39253 N39254 10
D39254 N39254 0 diode
R39255 N39254 N39255 10
D39255 N39255 0 diode
R39256 N39255 N39256 10
D39256 N39256 0 diode
R39257 N39256 N39257 10
D39257 N39257 0 diode
R39258 N39257 N39258 10
D39258 N39258 0 diode
R39259 N39258 N39259 10
D39259 N39259 0 diode
R39260 N39259 N39260 10
D39260 N39260 0 diode
R39261 N39260 N39261 10
D39261 N39261 0 diode
R39262 N39261 N39262 10
D39262 N39262 0 diode
R39263 N39262 N39263 10
D39263 N39263 0 diode
R39264 N39263 N39264 10
D39264 N39264 0 diode
R39265 N39264 N39265 10
D39265 N39265 0 diode
R39266 N39265 N39266 10
D39266 N39266 0 diode
R39267 N39266 N39267 10
D39267 N39267 0 diode
R39268 N39267 N39268 10
D39268 N39268 0 diode
R39269 N39268 N39269 10
D39269 N39269 0 diode
R39270 N39269 N39270 10
D39270 N39270 0 diode
R39271 N39270 N39271 10
D39271 N39271 0 diode
R39272 N39271 N39272 10
D39272 N39272 0 diode
R39273 N39272 N39273 10
D39273 N39273 0 diode
R39274 N39273 N39274 10
D39274 N39274 0 diode
R39275 N39274 N39275 10
D39275 N39275 0 diode
R39276 N39275 N39276 10
D39276 N39276 0 diode
R39277 N39276 N39277 10
D39277 N39277 0 diode
R39278 N39277 N39278 10
D39278 N39278 0 diode
R39279 N39278 N39279 10
D39279 N39279 0 diode
R39280 N39279 N39280 10
D39280 N39280 0 diode
R39281 N39280 N39281 10
D39281 N39281 0 diode
R39282 N39281 N39282 10
D39282 N39282 0 diode
R39283 N39282 N39283 10
D39283 N39283 0 diode
R39284 N39283 N39284 10
D39284 N39284 0 diode
R39285 N39284 N39285 10
D39285 N39285 0 diode
R39286 N39285 N39286 10
D39286 N39286 0 diode
R39287 N39286 N39287 10
D39287 N39287 0 diode
R39288 N39287 N39288 10
D39288 N39288 0 diode
R39289 N39288 N39289 10
D39289 N39289 0 diode
R39290 N39289 N39290 10
D39290 N39290 0 diode
R39291 N39290 N39291 10
D39291 N39291 0 diode
R39292 N39291 N39292 10
D39292 N39292 0 diode
R39293 N39292 N39293 10
D39293 N39293 0 diode
R39294 N39293 N39294 10
D39294 N39294 0 diode
R39295 N39294 N39295 10
D39295 N39295 0 diode
R39296 N39295 N39296 10
D39296 N39296 0 diode
R39297 N39296 N39297 10
D39297 N39297 0 diode
R39298 N39297 N39298 10
D39298 N39298 0 diode
R39299 N39298 N39299 10
D39299 N39299 0 diode
R39300 N39299 N39300 10
D39300 N39300 0 diode
R39301 N39300 N39301 10
D39301 N39301 0 diode
R39302 N39301 N39302 10
D39302 N39302 0 diode
R39303 N39302 N39303 10
D39303 N39303 0 diode
R39304 N39303 N39304 10
D39304 N39304 0 diode
R39305 N39304 N39305 10
D39305 N39305 0 diode
R39306 N39305 N39306 10
D39306 N39306 0 diode
R39307 N39306 N39307 10
D39307 N39307 0 diode
R39308 N39307 N39308 10
D39308 N39308 0 diode
R39309 N39308 N39309 10
D39309 N39309 0 diode
R39310 N39309 N39310 10
D39310 N39310 0 diode
R39311 N39310 N39311 10
D39311 N39311 0 diode
R39312 N39311 N39312 10
D39312 N39312 0 diode
R39313 N39312 N39313 10
D39313 N39313 0 diode
R39314 N39313 N39314 10
D39314 N39314 0 diode
R39315 N39314 N39315 10
D39315 N39315 0 diode
R39316 N39315 N39316 10
D39316 N39316 0 diode
R39317 N39316 N39317 10
D39317 N39317 0 diode
R39318 N39317 N39318 10
D39318 N39318 0 diode
R39319 N39318 N39319 10
D39319 N39319 0 diode
R39320 N39319 N39320 10
D39320 N39320 0 diode
R39321 N39320 N39321 10
D39321 N39321 0 diode
R39322 N39321 N39322 10
D39322 N39322 0 diode
R39323 N39322 N39323 10
D39323 N39323 0 diode
R39324 N39323 N39324 10
D39324 N39324 0 diode
R39325 N39324 N39325 10
D39325 N39325 0 diode
R39326 N39325 N39326 10
D39326 N39326 0 diode
R39327 N39326 N39327 10
D39327 N39327 0 diode
R39328 N39327 N39328 10
D39328 N39328 0 diode
R39329 N39328 N39329 10
D39329 N39329 0 diode
R39330 N39329 N39330 10
D39330 N39330 0 diode
R39331 N39330 N39331 10
D39331 N39331 0 diode
R39332 N39331 N39332 10
D39332 N39332 0 diode
R39333 N39332 N39333 10
D39333 N39333 0 diode
R39334 N39333 N39334 10
D39334 N39334 0 diode
R39335 N39334 N39335 10
D39335 N39335 0 diode
R39336 N39335 N39336 10
D39336 N39336 0 diode
R39337 N39336 N39337 10
D39337 N39337 0 diode
R39338 N39337 N39338 10
D39338 N39338 0 diode
R39339 N39338 N39339 10
D39339 N39339 0 diode
R39340 N39339 N39340 10
D39340 N39340 0 diode
R39341 N39340 N39341 10
D39341 N39341 0 diode
R39342 N39341 N39342 10
D39342 N39342 0 diode
R39343 N39342 N39343 10
D39343 N39343 0 diode
R39344 N39343 N39344 10
D39344 N39344 0 diode
R39345 N39344 N39345 10
D39345 N39345 0 diode
R39346 N39345 N39346 10
D39346 N39346 0 diode
R39347 N39346 N39347 10
D39347 N39347 0 diode
R39348 N39347 N39348 10
D39348 N39348 0 diode
R39349 N39348 N39349 10
D39349 N39349 0 diode
R39350 N39349 N39350 10
D39350 N39350 0 diode
R39351 N39350 N39351 10
D39351 N39351 0 diode
R39352 N39351 N39352 10
D39352 N39352 0 diode
R39353 N39352 N39353 10
D39353 N39353 0 diode
R39354 N39353 N39354 10
D39354 N39354 0 diode
R39355 N39354 N39355 10
D39355 N39355 0 diode
R39356 N39355 N39356 10
D39356 N39356 0 diode
R39357 N39356 N39357 10
D39357 N39357 0 diode
R39358 N39357 N39358 10
D39358 N39358 0 diode
R39359 N39358 N39359 10
D39359 N39359 0 diode
R39360 N39359 N39360 10
D39360 N39360 0 diode
R39361 N39360 N39361 10
D39361 N39361 0 diode
R39362 N39361 N39362 10
D39362 N39362 0 diode
R39363 N39362 N39363 10
D39363 N39363 0 diode
R39364 N39363 N39364 10
D39364 N39364 0 diode
R39365 N39364 N39365 10
D39365 N39365 0 diode
R39366 N39365 N39366 10
D39366 N39366 0 diode
R39367 N39366 N39367 10
D39367 N39367 0 diode
R39368 N39367 N39368 10
D39368 N39368 0 diode
R39369 N39368 N39369 10
D39369 N39369 0 diode
R39370 N39369 N39370 10
D39370 N39370 0 diode
R39371 N39370 N39371 10
D39371 N39371 0 diode
R39372 N39371 N39372 10
D39372 N39372 0 diode
R39373 N39372 N39373 10
D39373 N39373 0 diode
R39374 N39373 N39374 10
D39374 N39374 0 diode
R39375 N39374 N39375 10
D39375 N39375 0 diode
R39376 N39375 N39376 10
D39376 N39376 0 diode
R39377 N39376 N39377 10
D39377 N39377 0 diode
R39378 N39377 N39378 10
D39378 N39378 0 diode
R39379 N39378 N39379 10
D39379 N39379 0 diode
R39380 N39379 N39380 10
D39380 N39380 0 diode
R39381 N39380 N39381 10
D39381 N39381 0 diode
R39382 N39381 N39382 10
D39382 N39382 0 diode
R39383 N39382 N39383 10
D39383 N39383 0 diode
R39384 N39383 N39384 10
D39384 N39384 0 diode
R39385 N39384 N39385 10
D39385 N39385 0 diode
R39386 N39385 N39386 10
D39386 N39386 0 diode
R39387 N39386 N39387 10
D39387 N39387 0 diode
R39388 N39387 N39388 10
D39388 N39388 0 diode
R39389 N39388 N39389 10
D39389 N39389 0 diode
R39390 N39389 N39390 10
D39390 N39390 0 diode
R39391 N39390 N39391 10
D39391 N39391 0 diode
R39392 N39391 N39392 10
D39392 N39392 0 diode
R39393 N39392 N39393 10
D39393 N39393 0 diode
R39394 N39393 N39394 10
D39394 N39394 0 diode
R39395 N39394 N39395 10
D39395 N39395 0 diode
R39396 N39395 N39396 10
D39396 N39396 0 diode
R39397 N39396 N39397 10
D39397 N39397 0 diode
R39398 N39397 N39398 10
D39398 N39398 0 diode
R39399 N39398 N39399 10
D39399 N39399 0 diode
R39400 N39399 N39400 10
D39400 N39400 0 diode
R39401 N39400 N39401 10
D39401 N39401 0 diode
R39402 N39401 N39402 10
D39402 N39402 0 diode
R39403 N39402 N39403 10
D39403 N39403 0 diode
R39404 N39403 N39404 10
D39404 N39404 0 diode
R39405 N39404 N39405 10
D39405 N39405 0 diode
R39406 N39405 N39406 10
D39406 N39406 0 diode
R39407 N39406 N39407 10
D39407 N39407 0 diode
R39408 N39407 N39408 10
D39408 N39408 0 diode
R39409 N39408 N39409 10
D39409 N39409 0 diode
R39410 N39409 N39410 10
D39410 N39410 0 diode
R39411 N39410 N39411 10
D39411 N39411 0 diode
R39412 N39411 N39412 10
D39412 N39412 0 diode
R39413 N39412 N39413 10
D39413 N39413 0 diode
R39414 N39413 N39414 10
D39414 N39414 0 diode
R39415 N39414 N39415 10
D39415 N39415 0 diode
R39416 N39415 N39416 10
D39416 N39416 0 diode
R39417 N39416 N39417 10
D39417 N39417 0 diode
R39418 N39417 N39418 10
D39418 N39418 0 diode
R39419 N39418 N39419 10
D39419 N39419 0 diode
R39420 N39419 N39420 10
D39420 N39420 0 diode
R39421 N39420 N39421 10
D39421 N39421 0 diode
R39422 N39421 N39422 10
D39422 N39422 0 diode
R39423 N39422 N39423 10
D39423 N39423 0 diode
R39424 N39423 N39424 10
D39424 N39424 0 diode
R39425 N39424 N39425 10
D39425 N39425 0 diode
R39426 N39425 N39426 10
D39426 N39426 0 diode
R39427 N39426 N39427 10
D39427 N39427 0 diode
R39428 N39427 N39428 10
D39428 N39428 0 diode
R39429 N39428 N39429 10
D39429 N39429 0 diode
R39430 N39429 N39430 10
D39430 N39430 0 diode
R39431 N39430 N39431 10
D39431 N39431 0 diode
R39432 N39431 N39432 10
D39432 N39432 0 diode
R39433 N39432 N39433 10
D39433 N39433 0 diode
R39434 N39433 N39434 10
D39434 N39434 0 diode
R39435 N39434 N39435 10
D39435 N39435 0 diode
R39436 N39435 N39436 10
D39436 N39436 0 diode
R39437 N39436 N39437 10
D39437 N39437 0 diode
R39438 N39437 N39438 10
D39438 N39438 0 diode
R39439 N39438 N39439 10
D39439 N39439 0 diode
R39440 N39439 N39440 10
D39440 N39440 0 diode
R39441 N39440 N39441 10
D39441 N39441 0 diode
R39442 N39441 N39442 10
D39442 N39442 0 diode
R39443 N39442 N39443 10
D39443 N39443 0 diode
R39444 N39443 N39444 10
D39444 N39444 0 diode
R39445 N39444 N39445 10
D39445 N39445 0 diode
R39446 N39445 N39446 10
D39446 N39446 0 diode
R39447 N39446 N39447 10
D39447 N39447 0 diode
R39448 N39447 N39448 10
D39448 N39448 0 diode
R39449 N39448 N39449 10
D39449 N39449 0 diode
R39450 N39449 N39450 10
D39450 N39450 0 diode
R39451 N39450 N39451 10
D39451 N39451 0 diode
R39452 N39451 N39452 10
D39452 N39452 0 diode
R39453 N39452 N39453 10
D39453 N39453 0 diode
R39454 N39453 N39454 10
D39454 N39454 0 diode
R39455 N39454 N39455 10
D39455 N39455 0 diode
R39456 N39455 N39456 10
D39456 N39456 0 diode
R39457 N39456 N39457 10
D39457 N39457 0 diode
R39458 N39457 N39458 10
D39458 N39458 0 diode
R39459 N39458 N39459 10
D39459 N39459 0 diode
R39460 N39459 N39460 10
D39460 N39460 0 diode
R39461 N39460 N39461 10
D39461 N39461 0 diode
R39462 N39461 N39462 10
D39462 N39462 0 diode
R39463 N39462 N39463 10
D39463 N39463 0 diode
R39464 N39463 N39464 10
D39464 N39464 0 diode
R39465 N39464 N39465 10
D39465 N39465 0 diode
R39466 N39465 N39466 10
D39466 N39466 0 diode
R39467 N39466 N39467 10
D39467 N39467 0 diode
R39468 N39467 N39468 10
D39468 N39468 0 diode
R39469 N39468 N39469 10
D39469 N39469 0 diode
R39470 N39469 N39470 10
D39470 N39470 0 diode
R39471 N39470 N39471 10
D39471 N39471 0 diode
R39472 N39471 N39472 10
D39472 N39472 0 diode
R39473 N39472 N39473 10
D39473 N39473 0 diode
R39474 N39473 N39474 10
D39474 N39474 0 diode
R39475 N39474 N39475 10
D39475 N39475 0 diode
R39476 N39475 N39476 10
D39476 N39476 0 diode
R39477 N39476 N39477 10
D39477 N39477 0 diode
R39478 N39477 N39478 10
D39478 N39478 0 diode
R39479 N39478 N39479 10
D39479 N39479 0 diode
R39480 N39479 N39480 10
D39480 N39480 0 diode
R39481 N39480 N39481 10
D39481 N39481 0 diode
R39482 N39481 N39482 10
D39482 N39482 0 diode
R39483 N39482 N39483 10
D39483 N39483 0 diode
R39484 N39483 N39484 10
D39484 N39484 0 diode
R39485 N39484 N39485 10
D39485 N39485 0 diode
R39486 N39485 N39486 10
D39486 N39486 0 diode
R39487 N39486 N39487 10
D39487 N39487 0 diode
R39488 N39487 N39488 10
D39488 N39488 0 diode
R39489 N39488 N39489 10
D39489 N39489 0 diode
R39490 N39489 N39490 10
D39490 N39490 0 diode
R39491 N39490 N39491 10
D39491 N39491 0 diode
R39492 N39491 N39492 10
D39492 N39492 0 diode
R39493 N39492 N39493 10
D39493 N39493 0 diode
R39494 N39493 N39494 10
D39494 N39494 0 diode
R39495 N39494 N39495 10
D39495 N39495 0 diode
R39496 N39495 N39496 10
D39496 N39496 0 diode
R39497 N39496 N39497 10
D39497 N39497 0 diode
R39498 N39497 N39498 10
D39498 N39498 0 diode
R39499 N39498 N39499 10
D39499 N39499 0 diode
R39500 N39499 N39500 10
D39500 N39500 0 diode
R39501 N39500 N39501 10
D39501 N39501 0 diode
R39502 N39501 N39502 10
D39502 N39502 0 diode
R39503 N39502 N39503 10
D39503 N39503 0 diode
R39504 N39503 N39504 10
D39504 N39504 0 diode
R39505 N39504 N39505 10
D39505 N39505 0 diode
R39506 N39505 N39506 10
D39506 N39506 0 diode
R39507 N39506 N39507 10
D39507 N39507 0 diode
R39508 N39507 N39508 10
D39508 N39508 0 diode
R39509 N39508 N39509 10
D39509 N39509 0 diode
R39510 N39509 N39510 10
D39510 N39510 0 diode
R39511 N39510 N39511 10
D39511 N39511 0 diode
R39512 N39511 N39512 10
D39512 N39512 0 diode
R39513 N39512 N39513 10
D39513 N39513 0 diode
R39514 N39513 N39514 10
D39514 N39514 0 diode
R39515 N39514 N39515 10
D39515 N39515 0 diode
R39516 N39515 N39516 10
D39516 N39516 0 diode
R39517 N39516 N39517 10
D39517 N39517 0 diode
R39518 N39517 N39518 10
D39518 N39518 0 diode
R39519 N39518 N39519 10
D39519 N39519 0 diode
R39520 N39519 N39520 10
D39520 N39520 0 diode
R39521 N39520 N39521 10
D39521 N39521 0 diode
R39522 N39521 N39522 10
D39522 N39522 0 diode
R39523 N39522 N39523 10
D39523 N39523 0 diode
R39524 N39523 N39524 10
D39524 N39524 0 diode
R39525 N39524 N39525 10
D39525 N39525 0 diode
R39526 N39525 N39526 10
D39526 N39526 0 diode
R39527 N39526 N39527 10
D39527 N39527 0 diode
R39528 N39527 N39528 10
D39528 N39528 0 diode
R39529 N39528 N39529 10
D39529 N39529 0 diode
R39530 N39529 N39530 10
D39530 N39530 0 diode
R39531 N39530 N39531 10
D39531 N39531 0 diode
R39532 N39531 N39532 10
D39532 N39532 0 diode
R39533 N39532 N39533 10
D39533 N39533 0 diode
R39534 N39533 N39534 10
D39534 N39534 0 diode
R39535 N39534 N39535 10
D39535 N39535 0 diode
R39536 N39535 N39536 10
D39536 N39536 0 diode
R39537 N39536 N39537 10
D39537 N39537 0 diode
R39538 N39537 N39538 10
D39538 N39538 0 diode
R39539 N39538 N39539 10
D39539 N39539 0 diode
R39540 N39539 N39540 10
D39540 N39540 0 diode
R39541 N39540 N39541 10
D39541 N39541 0 diode
R39542 N39541 N39542 10
D39542 N39542 0 diode
R39543 N39542 N39543 10
D39543 N39543 0 diode
R39544 N39543 N39544 10
D39544 N39544 0 diode
R39545 N39544 N39545 10
D39545 N39545 0 diode
R39546 N39545 N39546 10
D39546 N39546 0 diode
R39547 N39546 N39547 10
D39547 N39547 0 diode
R39548 N39547 N39548 10
D39548 N39548 0 diode
R39549 N39548 N39549 10
D39549 N39549 0 diode
R39550 N39549 N39550 10
D39550 N39550 0 diode
R39551 N39550 N39551 10
D39551 N39551 0 diode
R39552 N39551 N39552 10
D39552 N39552 0 diode
R39553 N39552 N39553 10
D39553 N39553 0 diode
R39554 N39553 N39554 10
D39554 N39554 0 diode
R39555 N39554 N39555 10
D39555 N39555 0 diode
R39556 N39555 N39556 10
D39556 N39556 0 diode
R39557 N39556 N39557 10
D39557 N39557 0 diode
R39558 N39557 N39558 10
D39558 N39558 0 diode
R39559 N39558 N39559 10
D39559 N39559 0 diode
R39560 N39559 N39560 10
D39560 N39560 0 diode
R39561 N39560 N39561 10
D39561 N39561 0 diode
R39562 N39561 N39562 10
D39562 N39562 0 diode
R39563 N39562 N39563 10
D39563 N39563 0 diode
R39564 N39563 N39564 10
D39564 N39564 0 diode
R39565 N39564 N39565 10
D39565 N39565 0 diode
R39566 N39565 N39566 10
D39566 N39566 0 diode
R39567 N39566 N39567 10
D39567 N39567 0 diode
R39568 N39567 N39568 10
D39568 N39568 0 diode
R39569 N39568 N39569 10
D39569 N39569 0 diode
R39570 N39569 N39570 10
D39570 N39570 0 diode
R39571 N39570 N39571 10
D39571 N39571 0 diode
R39572 N39571 N39572 10
D39572 N39572 0 diode
R39573 N39572 N39573 10
D39573 N39573 0 diode
R39574 N39573 N39574 10
D39574 N39574 0 diode
R39575 N39574 N39575 10
D39575 N39575 0 diode
R39576 N39575 N39576 10
D39576 N39576 0 diode
R39577 N39576 N39577 10
D39577 N39577 0 diode
R39578 N39577 N39578 10
D39578 N39578 0 diode
R39579 N39578 N39579 10
D39579 N39579 0 diode
R39580 N39579 N39580 10
D39580 N39580 0 diode
R39581 N39580 N39581 10
D39581 N39581 0 diode
R39582 N39581 N39582 10
D39582 N39582 0 diode
R39583 N39582 N39583 10
D39583 N39583 0 diode
R39584 N39583 N39584 10
D39584 N39584 0 diode
R39585 N39584 N39585 10
D39585 N39585 0 diode
R39586 N39585 N39586 10
D39586 N39586 0 diode
R39587 N39586 N39587 10
D39587 N39587 0 diode
R39588 N39587 N39588 10
D39588 N39588 0 diode
R39589 N39588 N39589 10
D39589 N39589 0 diode
R39590 N39589 N39590 10
D39590 N39590 0 diode
R39591 N39590 N39591 10
D39591 N39591 0 diode
R39592 N39591 N39592 10
D39592 N39592 0 diode
R39593 N39592 N39593 10
D39593 N39593 0 diode
R39594 N39593 N39594 10
D39594 N39594 0 diode
R39595 N39594 N39595 10
D39595 N39595 0 diode
R39596 N39595 N39596 10
D39596 N39596 0 diode
R39597 N39596 N39597 10
D39597 N39597 0 diode
R39598 N39597 N39598 10
D39598 N39598 0 diode
R39599 N39598 N39599 10
D39599 N39599 0 diode
R39600 N39599 N39600 10
D39600 N39600 0 diode
R39601 N39600 N39601 10
D39601 N39601 0 diode
R39602 N39601 N39602 10
D39602 N39602 0 diode
R39603 N39602 N39603 10
D39603 N39603 0 diode
R39604 N39603 N39604 10
D39604 N39604 0 diode
R39605 N39604 N39605 10
D39605 N39605 0 diode
R39606 N39605 N39606 10
D39606 N39606 0 diode
R39607 N39606 N39607 10
D39607 N39607 0 diode
R39608 N39607 N39608 10
D39608 N39608 0 diode
R39609 N39608 N39609 10
D39609 N39609 0 diode
R39610 N39609 N39610 10
D39610 N39610 0 diode
R39611 N39610 N39611 10
D39611 N39611 0 diode
R39612 N39611 N39612 10
D39612 N39612 0 diode
R39613 N39612 N39613 10
D39613 N39613 0 diode
R39614 N39613 N39614 10
D39614 N39614 0 diode
R39615 N39614 N39615 10
D39615 N39615 0 diode
R39616 N39615 N39616 10
D39616 N39616 0 diode
R39617 N39616 N39617 10
D39617 N39617 0 diode
R39618 N39617 N39618 10
D39618 N39618 0 diode
R39619 N39618 N39619 10
D39619 N39619 0 diode
R39620 N39619 N39620 10
D39620 N39620 0 diode
R39621 N39620 N39621 10
D39621 N39621 0 diode
R39622 N39621 N39622 10
D39622 N39622 0 diode
R39623 N39622 N39623 10
D39623 N39623 0 diode
R39624 N39623 N39624 10
D39624 N39624 0 diode
R39625 N39624 N39625 10
D39625 N39625 0 diode
R39626 N39625 N39626 10
D39626 N39626 0 diode
R39627 N39626 N39627 10
D39627 N39627 0 diode
R39628 N39627 N39628 10
D39628 N39628 0 diode
R39629 N39628 N39629 10
D39629 N39629 0 diode
R39630 N39629 N39630 10
D39630 N39630 0 diode
R39631 N39630 N39631 10
D39631 N39631 0 diode
R39632 N39631 N39632 10
D39632 N39632 0 diode
R39633 N39632 N39633 10
D39633 N39633 0 diode
R39634 N39633 N39634 10
D39634 N39634 0 diode
R39635 N39634 N39635 10
D39635 N39635 0 diode
R39636 N39635 N39636 10
D39636 N39636 0 diode
R39637 N39636 N39637 10
D39637 N39637 0 diode
R39638 N39637 N39638 10
D39638 N39638 0 diode
R39639 N39638 N39639 10
D39639 N39639 0 diode
R39640 N39639 N39640 10
D39640 N39640 0 diode
R39641 N39640 N39641 10
D39641 N39641 0 diode
R39642 N39641 N39642 10
D39642 N39642 0 diode
R39643 N39642 N39643 10
D39643 N39643 0 diode
R39644 N39643 N39644 10
D39644 N39644 0 diode
R39645 N39644 N39645 10
D39645 N39645 0 diode
R39646 N39645 N39646 10
D39646 N39646 0 diode
R39647 N39646 N39647 10
D39647 N39647 0 diode
R39648 N39647 N39648 10
D39648 N39648 0 diode
R39649 N39648 N39649 10
D39649 N39649 0 diode
R39650 N39649 N39650 10
D39650 N39650 0 diode
R39651 N39650 N39651 10
D39651 N39651 0 diode
R39652 N39651 N39652 10
D39652 N39652 0 diode
R39653 N39652 N39653 10
D39653 N39653 0 diode
R39654 N39653 N39654 10
D39654 N39654 0 diode
R39655 N39654 N39655 10
D39655 N39655 0 diode
R39656 N39655 N39656 10
D39656 N39656 0 diode
R39657 N39656 N39657 10
D39657 N39657 0 diode
R39658 N39657 N39658 10
D39658 N39658 0 diode
R39659 N39658 N39659 10
D39659 N39659 0 diode
R39660 N39659 N39660 10
D39660 N39660 0 diode
R39661 N39660 N39661 10
D39661 N39661 0 diode
R39662 N39661 N39662 10
D39662 N39662 0 diode
R39663 N39662 N39663 10
D39663 N39663 0 diode
R39664 N39663 N39664 10
D39664 N39664 0 diode
R39665 N39664 N39665 10
D39665 N39665 0 diode
R39666 N39665 N39666 10
D39666 N39666 0 diode
R39667 N39666 N39667 10
D39667 N39667 0 diode
R39668 N39667 N39668 10
D39668 N39668 0 diode
R39669 N39668 N39669 10
D39669 N39669 0 diode
R39670 N39669 N39670 10
D39670 N39670 0 diode
R39671 N39670 N39671 10
D39671 N39671 0 diode
R39672 N39671 N39672 10
D39672 N39672 0 diode
R39673 N39672 N39673 10
D39673 N39673 0 diode
R39674 N39673 N39674 10
D39674 N39674 0 diode
R39675 N39674 N39675 10
D39675 N39675 0 diode
R39676 N39675 N39676 10
D39676 N39676 0 diode
R39677 N39676 N39677 10
D39677 N39677 0 diode
R39678 N39677 N39678 10
D39678 N39678 0 diode
R39679 N39678 N39679 10
D39679 N39679 0 diode
R39680 N39679 N39680 10
D39680 N39680 0 diode
R39681 N39680 N39681 10
D39681 N39681 0 diode
R39682 N39681 N39682 10
D39682 N39682 0 diode
R39683 N39682 N39683 10
D39683 N39683 0 diode
R39684 N39683 N39684 10
D39684 N39684 0 diode
R39685 N39684 N39685 10
D39685 N39685 0 diode
R39686 N39685 N39686 10
D39686 N39686 0 diode
R39687 N39686 N39687 10
D39687 N39687 0 diode
R39688 N39687 N39688 10
D39688 N39688 0 diode
R39689 N39688 N39689 10
D39689 N39689 0 diode
R39690 N39689 N39690 10
D39690 N39690 0 diode
R39691 N39690 N39691 10
D39691 N39691 0 diode
R39692 N39691 N39692 10
D39692 N39692 0 diode
R39693 N39692 N39693 10
D39693 N39693 0 diode
R39694 N39693 N39694 10
D39694 N39694 0 diode
R39695 N39694 N39695 10
D39695 N39695 0 diode
R39696 N39695 N39696 10
D39696 N39696 0 diode
R39697 N39696 N39697 10
D39697 N39697 0 diode
R39698 N39697 N39698 10
D39698 N39698 0 diode
R39699 N39698 N39699 10
D39699 N39699 0 diode
R39700 N39699 N39700 10
D39700 N39700 0 diode
R39701 N39700 N39701 10
D39701 N39701 0 diode
R39702 N39701 N39702 10
D39702 N39702 0 diode
R39703 N39702 N39703 10
D39703 N39703 0 diode
R39704 N39703 N39704 10
D39704 N39704 0 diode
R39705 N39704 N39705 10
D39705 N39705 0 diode
R39706 N39705 N39706 10
D39706 N39706 0 diode
R39707 N39706 N39707 10
D39707 N39707 0 diode
R39708 N39707 N39708 10
D39708 N39708 0 diode
R39709 N39708 N39709 10
D39709 N39709 0 diode
R39710 N39709 N39710 10
D39710 N39710 0 diode
R39711 N39710 N39711 10
D39711 N39711 0 diode
R39712 N39711 N39712 10
D39712 N39712 0 diode
R39713 N39712 N39713 10
D39713 N39713 0 diode
R39714 N39713 N39714 10
D39714 N39714 0 diode
R39715 N39714 N39715 10
D39715 N39715 0 diode
R39716 N39715 N39716 10
D39716 N39716 0 diode
R39717 N39716 N39717 10
D39717 N39717 0 diode
R39718 N39717 N39718 10
D39718 N39718 0 diode
R39719 N39718 N39719 10
D39719 N39719 0 diode
R39720 N39719 N39720 10
D39720 N39720 0 diode
R39721 N39720 N39721 10
D39721 N39721 0 diode
R39722 N39721 N39722 10
D39722 N39722 0 diode
R39723 N39722 N39723 10
D39723 N39723 0 diode
R39724 N39723 N39724 10
D39724 N39724 0 diode
R39725 N39724 N39725 10
D39725 N39725 0 diode
R39726 N39725 N39726 10
D39726 N39726 0 diode
R39727 N39726 N39727 10
D39727 N39727 0 diode
R39728 N39727 N39728 10
D39728 N39728 0 diode
R39729 N39728 N39729 10
D39729 N39729 0 diode
R39730 N39729 N39730 10
D39730 N39730 0 diode
R39731 N39730 N39731 10
D39731 N39731 0 diode
R39732 N39731 N39732 10
D39732 N39732 0 diode
R39733 N39732 N39733 10
D39733 N39733 0 diode
R39734 N39733 N39734 10
D39734 N39734 0 diode
R39735 N39734 N39735 10
D39735 N39735 0 diode
R39736 N39735 N39736 10
D39736 N39736 0 diode
R39737 N39736 N39737 10
D39737 N39737 0 diode
R39738 N39737 N39738 10
D39738 N39738 0 diode
R39739 N39738 N39739 10
D39739 N39739 0 diode
R39740 N39739 N39740 10
D39740 N39740 0 diode
R39741 N39740 N39741 10
D39741 N39741 0 diode
R39742 N39741 N39742 10
D39742 N39742 0 diode
R39743 N39742 N39743 10
D39743 N39743 0 diode
R39744 N39743 N39744 10
D39744 N39744 0 diode
R39745 N39744 N39745 10
D39745 N39745 0 diode
R39746 N39745 N39746 10
D39746 N39746 0 diode
R39747 N39746 N39747 10
D39747 N39747 0 diode
R39748 N39747 N39748 10
D39748 N39748 0 diode
R39749 N39748 N39749 10
D39749 N39749 0 diode
R39750 N39749 N39750 10
D39750 N39750 0 diode
R39751 N39750 N39751 10
D39751 N39751 0 diode
R39752 N39751 N39752 10
D39752 N39752 0 diode
R39753 N39752 N39753 10
D39753 N39753 0 diode
R39754 N39753 N39754 10
D39754 N39754 0 diode
R39755 N39754 N39755 10
D39755 N39755 0 diode
R39756 N39755 N39756 10
D39756 N39756 0 diode
R39757 N39756 N39757 10
D39757 N39757 0 diode
R39758 N39757 N39758 10
D39758 N39758 0 diode
R39759 N39758 N39759 10
D39759 N39759 0 diode
R39760 N39759 N39760 10
D39760 N39760 0 diode
R39761 N39760 N39761 10
D39761 N39761 0 diode
R39762 N39761 N39762 10
D39762 N39762 0 diode
R39763 N39762 N39763 10
D39763 N39763 0 diode
R39764 N39763 N39764 10
D39764 N39764 0 diode
R39765 N39764 N39765 10
D39765 N39765 0 diode
R39766 N39765 N39766 10
D39766 N39766 0 diode
R39767 N39766 N39767 10
D39767 N39767 0 diode
R39768 N39767 N39768 10
D39768 N39768 0 diode
R39769 N39768 N39769 10
D39769 N39769 0 diode
R39770 N39769 N39770 10
D39770 N39770 0 diode
R39771 N39770 N39771 10
D39771 N39771 0 diode
R39772 N39771 N39772 10
D39772 N39772 0 diode
R39773 N39772 N39773 10
D39773 N39773 0 diode
R39774 N39773 N39774 10
D39774 N39774 0 diode
R39775 N39774 N39775 10
D39775 N39775 0 diode
R39776 N39775 N39776 10
D39776 N39776 0 diode
R39777 N39776 N39777 10
D39777 N39777 0 diode
R39778 N39777 N39778 10
D39778 N39778 0 diode
R39779 N39778 N39779 10
D39779 N39779 0 diode
R39780 N39779 N39780 10
D39780 N39780 0 diode
R39781 N39780 N39781 10
D39781 N39781 0 diode
R39782 N39781 N39782 10
D39782 N39782 0 diode
R39783 N39782 N39783 10
D39783 N39783 0 diode
R39784 N39783 N39784 10
D39784 N39784 0 diode
R39785 N39784 N39785 10
D39785 N39785 0 diode
R39786 N39785 N39786 10
D39786 N39786 0 diode
R39787 N39786 N39787 10
D39787 N39787 0 diode
R39788 N39787 N39788 10
D39788 N39788 0 diode
R39789 N39788 N39789 10
D39789 N39789 0 diode
R39790 N39789 N39790 10
D39790 N39790 0 diode
R39791 N39790 N39791 10
D39791 N39791 0 diode
R39792 N39791 N39792 10
D39792 N39792 0 diode
R39793 N39792 N39793 10
D39793 N39793 0 diode
R39794 N39793 N39794 10
D39794 N39794 0 diode
R39795 N39794 N39795 10
D39795 N39795 0 diode
R39796 N39795 N39796 10
D39796 N39796 0 diode
R39797 N39796 N39797 10
D39797 N39797 0 diode
R39798 N39797 N39798 10
D39798 N39798 0 diode
R39799 N39798 N39799 10
D39799 N39799 0 diode
R39800 N39799 N39800 10
D39800 N39800 0 diode
R39801 N39800 N39801 10
D39801 N39801 0 diode
R39802 N39801 N39802 10
D39802 N39802 0 diode
R39803 N39802 N39803 10
D39803 N39803 0 diode
R39804 N39803 N39804 10
D39804 N39804 0 diode
R39805 N39804 N39805 10
D39805 N39805 0 diode
R39806 N39805 N39806 10
D39806 N39806 0 diode
R39807 N39806 N39807 10
D39807 N39807 0 diode
R39808 N39807 N39808 10
D39808 N39808 0 diode
R39809 N39808 N39809 10
D39809 N39809 0 diode
R39810 N39809 N39810 10
D39810 N39810 0 diode
R39811 N39810 N39811 10
D39811 N39811 0 diode
R39812 N39811 N39812 10
D39812 N39812 0 diode
R39813 N39812 N39813 10
D39813 N39813 0 diode
R39814 N39813 N39814 10
D39814 N39814 0 diode
R39815 N39814 N39815 10
D39815 N39815 0 diode
R39816 N39815 N39816 10
D39816 N39816 0 diode
R39817 N39816 N39817 10
D39817 N39817 0 diode
R39818 N39817 N39818 10
D39818 N39818 0 diode
R39819 N39818 N39819 10
D39819 N39819 0 diode
R39820 N39819 N39820 10
D39820 N39820 0 diode
R39821 N39820 N39821 10
D39821 N39821 0 diode
R39822 N39821 N39822 10
D39822 N39822 0 diode
R39823 N39822 N39823 10
D39823 N39823 0 diode
R39824 N39823 N39824 10
D39824 N39824 0 diode
R39825 N39824 N39825 10
D39825 N39825 0 diode
R39826 N39825 N39826 10
D39826 N39826 0 diode
R39827 N39826 N39827 10
D39827 N39827 0 diode
R39828 N39827 N39828 10
D39828 N39828 0 diode
R39829 N39828 N39829 10
D39829 N39829 0 diode
R39830 N39829 N39830 10
D39830 N39830 0 diode
R39831 N39830 N39831 10
D39831 N39831 0 diode
R39832 N39831 N39832 10
D39832 N39832 0 diode
R39833 N39832 N39833 10
D39833 N39833 0 diode
R39834 N39833 N39834 10
D39834 N39834 0 diode
R39835 N39834 N39835 10
D39835 N39835 0 diode
R39836 N39835 N39836 10
D39836 N39836 0 diode
R39837 N39836 N39837 10
D39837 N39837 0 diode
R39838 N39837 N39838 10
D39838 N39838 0 diode
R39839 N39838 N39839 10
D39839 N39839 0 diode
R39840 N39839 N39840 10
D39840 N39840 0 diode
R39841 N39840 N39841 10
D39841 N39841 0 diode
R39842 N39841 N39842 10
D39842 N39842 0 diode
R39843 N39842 N39843 10
D39843 N39843 0 diode
R39844 N39843 N39844 10
D39844 N39844 0 diode
R39845 N39844 N39845 10
D39845 N39845 0 diode
R39846 N39845 N39846 10
D39846 N39846 0 diode
R39847 N39846 N39847 10
D39847 N39847 0 diode
R39848 N39847 N39848 10
D39848 N39848 0 diode
R39849 N39848 N39849 10
D39849 N39849 0 diode
R39850 N39849 N39850 10
D39850 N39850 0 diode
R39851 N39850 N39851 10
D39851 N39851 0 diode
R39852 N39851 N39852 10
D39852 N39852 0 diode
R39853 N39852 N39853 10
D39853 N39853 0 diode
R39854 N39853 N39854 10
D39854 N39854 0 diode
R39855 N39854 N39855 10
D39855 N39855 0 diode
R39856 N39855 N39856 10
D39856 N39856 0 diode
R39857 N39856 N39857 10
D39857 N39857 0 diode
R39858 N39857 N39858 10
D39858 N39858 0 diode
R39859 N39858 N39859 10
D39859 N39859 0 diode
R39860 N39859 N39860 10
D39860 N39860 0 diode
R39861 N39860 N39861 10
D39861 N39861 0 diode
R39862 N39861 N39862 10
D39862 N39862 0 diode
R39863 N39862 N39863 10
D39863 N39863 0 diode
R39864 N39863 N39864 10
D39864 N39864 0 diode
R39865 N39864 N39865 10
D39865 N39865 0 diode
R39866 N39865 N39866 10
D39866 N39866 0 diode
R39867 N39866 N39867 10
D39867 N39867 0 diode
R39868 N39867 N39868 10
D39868 N39868 0 diode
R39869 N39868 N39869 10
D39869 N39869 0 diode
R39870 N39869 N39870 10
D39870 N39870 0 diode
R39871 N39870 N39871 10
D39871 N39871 0 diode
R39872 N39871 N39872 10
D39872 N39872 0 diode
R39873 N39872 N39873 10
D39873 N39873 0 diode
R39874 N39873 N39874 10
D39874 N39874 0 diode
R39875 N39874 N39875 10
D39875 N39875 0 diode
R39876 N39875 N39876 10
D39876 N39876 0 diode
R39877 N39876 N39877 10
D39877 N39877 0 diode
R39878 N39877 N39878 10
D39878 N39878 0 diode
R39879 N39878 N39879 10
D39879 N39879 0 diode
R39880 N39879 N39880 10
D39880 N39880 0 diode
R39881 N39880 N39881 10
D39881 N39881 0 diode
R39882 N39881 N39882 10
D39882 N39882 0 diode
R39883 N39882 N39883 10
D39883 N39883 0 diode
R39884 N39883 N39884 10
D39884 N39884 0 diode
R39885 N39884 N39885 10
D39885 N39885 0 diode
R39886 N39885 N39886 10
D39886 N39886 0 diode
R39887 N39886 N39887 10
D39887 N39887 0 diode
R39888 N39887 N39888 10
D39888 N39888 0 diode
R39889 N39888 N39889 10
D39889 N39889 0 diode
R39890 N39889 N39890 10
D39890 N39890 0 diode
R39891 N39890 N39891 10
D39891 N39891 0 diode
R39892 N39891 N39892 10
D39892 N39892 0 diode
R39893 N39892 N39893 10
D39893 N39893 0 diode
R39894 N39893 N39894 10
D39894 N39894 0 diode
R39895 N39894 N39895 10
D39895 N39895 0 diode
R39896 N39895 N39896 10
D39896 N39896 0 diode
R39897 N39896 N39897 10
D39897 N39897 0 diode
R39898 N39897 N39898 10
D39898 N39898 0 diode
R39899 N39898 N39899 10
D39899 N39899 0 diode
R39900 N39899 N39900 10
D39900 N39900 0 diode
R39901 N39900 N39901 10
D39901 N39901 0 diode
R39902 N39901 N39902 10
D39902 N39902 0 diode
R39903 N39902 N39903 10
D39903 N39903 0 diode
R39904 N39903 N39904 10
D39904 N39904 0 diode
R39905 N39904 N39905 10
D39905 N39905 0 diode
R39906 N39905 N39906 10
D39906 N39906 0 diode
R39907 N39906 N39907 10
D39907 N39907 0 diode
R39908 N39907 N39908 10
D39908 N39908 0 diode
R39909 N39908 N39909 10
D39909 N39909 0 diode
R39910 N39909 N39910 10
D39910 N39910 0 diode
R39911 N39910 N39911 10
D39911 N39911 0 diode
R39912 N39911 N39912 10
D39912 N39912 0 diode
R39913 N39912 N39913 10
D39913 N39913 0 diode
R39914 N39913 N39914 10
D39914 N39914 0 diode
R39915 N39914 N39915 10
D39915 N39915 0 diode
R39916 N39915 N39916 10
D39916 N39916 0 diode
R39917 N39916 N39917 10
D39917 N39917 0 diode
R39918 N39917 N39918 10
D39918 N39918 0 diode
R39919 N39918 N39919 10
D39919 N39919 0 diode
R39920 N39919 N39920 10
D39920 N39920 0 diode
R39921 N39920 N39921 10
D39921 N39921 0 diode
R39922 N39921 N39922 10
D39922 N39922 0 diode
R39923 N39922 N39923 10
D39923 N39923 0 diode
R39924 N39923 N39924 10
D39924 N39924 0 diode
R39925 N39924 N39925 10
D39925 N39925 0 diode
R39926 N39925 N39926 10
D39926 N39926 0 diode
R39927 N39926 N39927 10
D39927 N39927 0 diode
R39928 N39927 N39928 10
D39928 N39928 0 diode
R39929 N39928 N39929 10
D39929 N39929 0 diode
R39930 N39929 N39930 10
D39930 N39930 0 diode
R39931 N39930 N39931 10
D39931 N39931 0 diode
R39932 N39931 N39932 10
D39932 N39932 0 diode
R39933 N39932 N39933 10
D39933 N39933 0 diode
R39934 N39933 N39934 10
D39934 N39934 0 diode
R39935 N39934 N39935 10
D39935 N39935 0 diode
R39936 N39935 N39936 10
D39936 N39936 0 diode
R39937 N39936 N39937 10
D39937 N39937 0 diode
R39938 N39937 N39938 10
D39938 N39938 0 diode
R39939 N39938 N39939 10
D39939 N39939 0 diode
R39940 N39939 N39940 10
D39940 N39940 0 diode
R39941 N39940 N39941 10
D39941 N39941 0 diode
R39942 N39941 N39942 10
D39942 N39942 0 diode
R39943 N39942 N39943 10
D39943 N39943 0 diode
R39944 N39943 N39944 10
D39944 N39944 0 diode
R39945 N39944 N39945 10
D39945 N39945 0 diode
R39946 N39945 N39946 10
D39946 N39946 0 diode
R39947 N39946 N39947 10
D39947 N39947 0 diode
R39948 N39947 N39948 10
D39948 N39948 0 diode
R39949 N39948 N39949 10
D39949 N39949 0 diode
R39950 N39949 N39950 10
D39950 N39950 0 diode
R39951 N39950 N39951 10
D39951 N39951 0 diode
R39952 N39951 N39952 10
D39952 N39952 0 diode
R39953 N39952 N39953 10
D39953 N39953 0 diode
R39954 N39953 N39954 10
D39954 N39954 0 diode
R39955 N39954 N39955 10
D39955 N39955 0 diode
R39956 N39955 N39956 10
D39956 N39956 0 diode
R39957 N39956 N39957 10
D39957 N39957 0 diode
R39958 N39957 N39958 10
D39958 N39958 0 diode
R39959 N39958 N39959 10
D39959 N39959 0 diode
R39960 N39959 N39960 10
D39960 N39960 0 diode
R39961 N39960 N39961 10
D39961 N39961 0 diode
R39962 N39961 N39962 10
D39962 N39962 0 diode
R39963 N39962 N39963 10
D39963 N39963 0 diode
R39964 N39963 N39964 10
D39964 N39964 0 diode
R39965 N39964 N39965 10
D39965 N39965 0 diode
R39966 N39965 N39966 10
D39966 N39966 0 diode
R39967 N39966 N39967 10
D39967 N39967 0 diode
R39968 N39967 N39968 10
D39968 N39968 0 diode
R39969 N39968 N39969 10
D39969 N39969 0 diode
R39970 N39969 N39970 10
D39970 N39970 0 diode
R39971 N39970 N39971 10
D39971 N39971 0 diode
R39972 N39971 N39972 10
D39972 N39972 0 diode
R39973 N39972 N39973 10
D39973 N39973 0 diode
R39974 N39973 N39974 10
D39974 N39974 0 diode
R39975 N39974 N39975 10
D39975 N39975 0 diode
R39976 N39975 N39976 10
D39976 N39976 0 diode
R39977 N39976 N39977 10
D39977 N39977 0 diode
R39978 N39977 N39978 10
D39978 N39978 0 diode
R39979 N39978 N39979 10
D39979 N39979 0 diode
R39980 N39979 N39980 10
D39980 N39980 0 diode
R39981 N39980 N39981 10
D39981 N39981 0 diode
R39982 N39981 N39982 10
D39982 N39982 0 diode
R39983 N39982 N39983 10
D39983 N39983 0 diode
R39984 N39983 N39984 10
D39984 N39984 0 diode
R39985 N39984 N39985 10
D39985 N39985 0 diode
R39986 N39985 N39986 10
D39986 N39986 0 diode
R39987 N39986 N39987 10
D39987 N39987 0 diode
R39988 N39987 N39988 10
D39988 N39988 0 diode
R39989 N39988 N39989 10
D39989 N39989 0 diode
R39990 N39989 N39990 10
D39990 N39990 0 diode
R39991 N39990 N39991 10
D39991 N39991 0 diode
R39992 N39991 N39992 10
D39992 N39992 0 diode
R39993 N39992 N39993 10
D39993 N39993 0 diode
R39994 N39993 N39994 10
D39994 N39994 0 diode
R39995 N39994 N39995 10
D39995 N39995 0 diode
R39996 N39995 N39996 10
D39996 N39996 0 diode
R39997 N39996 N39997 10
D39997 N39997 0 diode
R39998 N39997 N39998 10
D39998 N39998 0 diode
R39999 N39998 N39999 10
D39999 N39999 0 diode
R40000 N39999 N40000 10
D40000 N40000 0 diode
R40001 N40000 N40001 10
D40001 N40001 0 diode
R40002 N40001 N40002 10
D40002 N40002 0 diode
R40003 N40002 N40003 10
D40003 N40003 0 diode
R40004 N40003 N40004 10
D40004 N40004 0 diode
R40005 N40004 N40005 10
D40005 N40005 0 diode
R40006 N40005 N40006 10
D40006 N40006 0 diode
R40007 N40006 N40007 10
D40007 N40007 0 diode
R40008 N40007 N40008 10
D40008 N40008 0 diode
R40009 N40008 N40009 10
D40009 N40009 0 diode
R40010 N40009 N40010 10
D40010 N40010 0 diode
R40011 N40010 N40011 10
D40011 N40011 0 diode
R40012 N40011 N40012 10
D40012 N40012 0 diode
R40013 N40012 N40013 10
D40013 N40013 0 diode
R40014 N40013 N40014 10
D40014 N40014 0 diode
R40015 N40014 N40015 10
D40015 N40015 0 diode
R40016 N40015 N40016 10
D40016 N40016 0 diode
R40017 N40016 N40017 10
D40017 N40017 0 diode
R40018 N40017 N40018 10
D40018 N40018 0 diode
R40019 N40018 N40019 10
D40019 N40019 0 diode
R40020 N40019 N40020 10
D40020 N40020 0 diode
R40021 N40020 N40021 10
D40021 N40021 0 diode
R40022 N40021 N40022 10
D40022 N40022 0 diode
R40023 N40022 N40023 10
D40023 N40023 0 diode
R40024 N40023 N40024 10
D40024 N40024 0 diode
R40025 N40024 N40025 10
D40025 N40025 0 diode
R40026 N40025 N40026 10
D40026 N40026 0 diode
R40027 N40026 N40027 10
D40027 N40027 0 diode
R40028 N40027 N40028 10
D40028 N40028 0 diode
R40029 N40028 N40029 10
D40029 N40029 0 diode
R40030 N40029 N40030 10
D40030 N40030 0 diode
R40031 N40030 N40031 10
D40031 N40031 0 diode
R40032 N40031 N40032 10
D40032 N40032 0 diode
R40033 N40032 N40033 10
D40033 N40033 0 diode
R40034 N40033 N40034 10
D40034 N40034 0 diode
R40035 N40034 N40035 10
D40035 N40035 0 diode
R40036 N40035 N40036 10
D40036 N40036 0 diode
R40037 N40036 N40037 10
D40037 N40037 0 diode
R40038 N40037 N40038 10
D40038 N40038 0 diode
R40039 N40038 N40039 10
D40039 N40039 0 diode
R40040 N40039 N40040 10
D40040 N40040 0 diode
R40041 N40040 N40041 10
D40041 N40041 0 diode
R40042 N40041 N40042 10
D40042 N40042 0 diode
R40043 N40042 N40043 10
D40043 N40043 0 diode
R40044 N40043 N40044 10
D40044 N40044 0 diode
R40045 N40044 N40045 10
D40045 N40045 0 diode
R40046 N40045 N40046 10
D40046 N40046 0 diode
R40047 N40046 N40047 10
D40047 N40047 0 diode
R40048 N40047 N40048 10
D40048 N40048 0 diode
R40049 N40048 N40049 10
D40049 N40049 0 diode
R40050 N40049 N40050 10
D40050 N40050 0 diode
R40051 N40050 N40051 10
D40051 N40051 0 diode
R40052 N40051 N40052 10
D40052 N40052 0 diode
R40053 N40052 N40053 10
D40053 N40053 0 diode
R40054 N40053 N40054 10
D40054 N40054 0 diode
R40055 N40054 N40055 10
D40055 N40055 0 diode
R40056 N40055 N40056 10
D40056 N40056 0 diode
R40057 N40056 N40057 10
D40057 N40057 0 diode
R40058 N40057 N40058 10
D40058 N40058 0 diode
R40059 N40058 N40059 10
D40059 N40059 0 diode
R40060 N40059 N40060 10
D40060 N40060 0 diode
R40061 N40060 N40061 10
D40061 N40061 0 diode
R40062 N40061 N40062 10
D40062 N40062 0 diode
R40063 N40062 N40063 10
D40063 N40063 0 diode
R40064 N40063 N40064 10
D40064 N40064 0 diode
R40065 N40064 N40065 10
D40065 N40065 0 diode
R40066 N40065 N40066 10
D40066 N40066 0 diode
R40067 N40066 N40067 10
D40067 N40067 0 diode
R40068 N40067 N40068 10
D40068 N40068 0 diode
R40069 N40068 N40069 10
D40069 N40069 0 diode
R40070 N40069 N40070 10
D40070 N40070 0 diode
R40071 N40070 N40071 10
D40071 N40071 0 diode
R40072 N40071 N40072 10
D40072 N40072 0 diode
R40073 N40072 N40073 10
D40073 N40073 0 diode
R40074 N40073 N40074 10
D40074 N40074 0 diode
R40075 N40074 N40075 10
D40075 N40075 0 diode
R40076 N40075 N40076 10
D40076 N40076 0 diode
R40077 N40076 N40077 10
D40077 N40077 0 diode
R40078 N40077 N40078 10
D40078 N40078 0 diode
R40079 N40078 N40079 10
D40079 N40079 0 diode
R40080 N40079 N40080 10
D40080 N40080 0 diode
R40081 N40080 N40081 10
D40081 N40081 0 diode
R40082 N40081 N40082 10
D40082 N40082 0 diode
R40083 N40082 N40083 10
D40083 N40083 0 diode
R40084 N40083 N40084 10
D40084 N40084 0 diode
R40085 N40084 N40085 10
D40085 N40085 0 diode
R40086 N40085 N40086 10
D40086 N40086 0 diode
R40087 N40086 N40087 10
D40087 N40087 0 diode
R40088 N40087 N40088 10
D40088 N40088 0 diode
R40089 N40088 N40089 10
D40089 N40089 0 diode
R40090 N40089 N40090 10
D40090 N40090 0 diode
R40091 N40090 N40091 10
D40091 N40091 0 diode
R40092 N40091 N40092 10
D40092 N40092 0 diode
R40093 N40092 N40093 10
D40093 N40093 0 diode
R40094 N40093 N40094 10
D40094 N40094 0 diode
R40095 N40094 N40095 10
D40095 N40095 0 diode
R40096 N40095 N40096 10
D40096 N40096 0 diode
R40097 N40096 N40097 10
D40097 N40097 0 diode
R40098 N40097 N40098 10
D40098 N40098 0 diode
R40099 N40098 N40099 10
D40099 N40099 0 diode
R40100 N40099 N40100 10
D40100 N40100 0 diode
R40101 N40100 N40101 10
D40101 N40101 0 diode
R40102 N40101 N40102 10
D40102 N40102 0 diode
R40103 N40102 N40103 10
D40103 N40103 0 diode
R40104 N40103 N40104 10
D40104 N40104 0 diode
R40105 N40104 N40105 10
D40105 N40105 0 diode
R40106 N40105 N40106 10
D40106 N40106 0 diode
R40107 N40106 N40107 10
D40107 N40107 0 diode
R40108 N40107 N40108 10
D40108 N40108 0 diode
R40109 N40108 N40109 10
D40109 N40109 0 diode
R40110 N40109 N40110 10
D40110 N40110 0 diode
R40111 N40110 N40111 10
D40111 N40111 0 diode
R40112 N40111 N40112 10
D40112 N40112 0 diode
R40113 N40112 N40113 10
D40113 N40113 0 diode
R40114 N40113 N40114 10
D40114 N40114 0 diode
R40115 N40114 N40115 10
D40115 N40115 0 diode
R40116 N40115 N40116 10
D40116 N40116 0 diode
R40117 N40116 N40117 10
D40117 N40117 0 diode
R40118 N40117 N40118 10
D40118 N40118 0 diode
R40119 N40118 N40119 10
D40119 N40119 0 diode
R40120 N40119 N40120 10
D40120 N40120 0 diode
R40121 N40120 N40121 10
D40121 N40121 0 diode
R40122 N40121 N40122 10
D40122 N40122 0 diode
R40123 N40122 N40123 10
D40123 N40123 0 diode
R40124 N40123 N40124 10
D40124 N40124 0 diode
R40125 N40124 N40125 10
D40125 N40125 0 diode
R40126 N40125 N40126 10
D40126 N40126 0 diode
R40127 N40126 N40127 10
D40127 N40127 0 diode
R40128 N40127 N40128 10
D40128 N40128 0 diode
R40129 N40128 N40129 10
D40129 N40129 0 diode
R40130 N40129 N40130 10
D40130 N40130 0 diode
R40131 N40130 N40131 10
D40131 N40131 0 diode
R40132 N40131 N40132 10
D40132 N40132 0 diode
R40133 N40132 N40133 10
D40133 N40133 0 diode
R40134 N40133 N40134 10
D40134 N40134 0 diode
R40135 N40134 N40135 10
D40135 N40135 0 diode
R40136 N40135 N40136 10
D40136 N40136 0 diode
R40137 N40136 N40137 10
D40137 N40137 0 diode
R40138 N40137 N40138 10
D40138 N40138 0 diode
R40139 N40138 N40139 10
D40139 N40139 0 diode
R40140 N40139 N40140 10
D40140 N40140 0 diode
R40141 N40140 N40141 10
D40141 N40141 0 diode
R40142 N40141 N40142 10
D40142 N40142 0 diode
R40143 N40142 N40143 10
D40143 N40143 0 diode
R40144 N40143 N40144 10
D40144 N40144 0 diode
R40145 N40144 N40145 10
D40145 N40145 0 diode
R40146 N40145 N40146 10
D40146 N40146 0 diode
R40147 N40146 N40147 10
D40147 N40147 0 diode
R40148 N40147 N40148 10
D40148 N40148 0 diode
R40149 N40148 N40149 10
D40149 N40149 0 diode
R40150 N40149 N40150 10
D40150 N40150 0 diode
R40151 N40150 N40151 10
D40151 N40151 0 diode
R40152 N40151 N40152 10
D40152 N40152 0 diode
R40153 N40152 N40153 10
D40153 N40153 0 diode
R40154 N40153 N40154 10
D40154 N40154 0 diode
R40155 N40154 N40155 10
D40155 N40155 0 diode
R40156 N40155 N40156 10
D40156 N40156 0 diode
R40157 N40156 N40157 10
D40157 N40157 0 diode
R40158 N40157 N40158 10
D40158 N40158 0 diode
R40159 N40158 N40159 10
D40159 N40159 0 diode
R40160 N40159 N40160 10
D40160 N40160 0 diode
R40161 N40160 N40161 10
D40161 N40161 0 diode
R40162 N40161 N40162 10
D40162 N40162 0 diode
R40163 N40162 N40163 10
D40163 N40163 0 diode
R40164 N40163 N40164 10
D40164 N40164 0 diode
R40165 N40164 N40165 10
D40165 N40165 0 diode
R40166 N40165 N40166 10
D40166 N40166 0 diode
R40167 N40166 N40167 10
D40167 N40167 0 diode
R40168 N40167 N40168 10
D40168 N40168 0 diode
R40169 N40168 N40169 10
D40169 N40169 0 diode
R40170 N40169 N40170 10
D40170 N40170 0 diode
R40171 N40170 N40171 10
D40171 N40171 0 diode
R40172 N40171 N40172 10
D40172 N40172 0 diode
R40173 N40172 N40173 10
D40173 N40173 0 diode
R40174 N40173 N40174 10
D40174 N40174 0 diode
R40175 N40174 N40175 10
D40175 N40175 0 diode
R40176 N40175 N40176 10
D40176 N40176 0 diode
R40177 N40176 N40177 10
D40177 N40177 0 diode
R40178 N40177 N40178 10
D40178 N40178 0 diode
R40179 N40178 N40179 10
D40179 N40179 0 diode
R40180 N40179 N40180 10
D40180 N40180 0 diode
R40181 N40180 N40181 10
D40181 N40181 0 diode
R40182 N40181 N40182 10
D40182 N40182 0 diode
R40183 N40182 N40183 10
D40183 N40183 0 diode
R40184 N40183 N40184 10
D40184 N40184 0 diode
R40185 N40184 N40185 10
D40185 N40185 0 diode
R40186 N40185 N40186 10
D40186 N40186 0 diode
R40187 N40186 N40187 10
D40187 N40187 0 diode
R40188 N40187 N40188 10
D40188 N40188 0 diode
R40189 N40188 N40189 10
D40189 N40189 0 diode
R40190 N40189 N40190 10
D40190 N40190 0 diode
R40191 N40190 N40191 10
D40191 N40191 0 diode
R40192 N40191 N40192 10
D40192 N40192 0 diode
R40193 N40192 N40193 10
D40193 N40193 0 diode
R40194 N40193 N40194 10
D40194 N40194 0 diode
R40195 N40194 N40195 10
D40195 N40195 0 diode
R40196 N40195 N40196 10
D40196 N40196 0 diode
R40197 N40196 N40197 10
D40197 N40197 0 diode
R40198 N40197 N40198 10
D40198 N40198 0 diode
R40199 N40198 N40199 10
D40199 N40199 0 diode
R40200 N40199 N40200 10
D40200 N40200 0 diode
R40201 N40200 N40201 10
D40201 N40201 0 diode
R40202 N40201 N40202 10
D40202 N40202 0 diode
R40203 N40202 N40203 10
D40203 N40203 0 diode
R40204 N40203 N40204 10
D40204 N40204 0 diode
R40205 N40204 N40205 10
D40205 N40205 0 diode
R40206 N40205 N40206 10
D40206 N40206 0 diode
R40207 N40206 N40207 10
D40207 N40207 0 diode
R40208 N40207 N40208 10
D40208 N40208 0 diode
R40209 N40208 N40209 10
D40209 N40209 0 diode
R40210 N40209 N40210 10
D40210 N40210 0 diode
R40211 N40210 N40211 10
D40211 N40211 0 diode
R40212 N40211 N40212 10
D40212 N40212 0 diode
R40213 N40212 N40213 10
D40213 N40213 0 diode
R40214 N40213 N40214 10
D40214 N40214 0 diode
R40215 N40214 N40215 10
D40215 N40215 0 diode
R40216 N40215 N40216 10
D40216 N40216 0 diode
R40217 N40216 N40217 10
D40217 N40217 0 diode
R40218 N40217 N40218 10
D40218 N40218 0 diode
R40219 N40218 N40219 10
D40219 N40219 0 diode
R40220 N40219 N40220 10
D40220 N40220 0 diode
R40221 N40220 N40221 10
D40221 N40221 0 diode
R40222 N40221 N40222 10
D40222 N40222 0 diode
R40223 N40222 N40223 10
D40223 N40223 0 diode
R40224 N40223 N40224 10
D40224 N40224 0 diode
R40225 N40224 N40225 10
D40225 N40225 0 diode
R40226 N40225 N40226 10
D40226 N40226 0 diode
R40227 N40226 N40227 10
D40227 N40227 0 diode
R40228 N40227 N40228 10
D40228 N40228 0 diode
R40229 N40228 N40229 10
D40229 N40229 0 diode
R40230 N40229 N40230 10
D40230 N40230 0 diode
R40231 N40230 N40231 10
D40231 N40231 0 diode
R40232 N40231 N40232 10
D40232 N40232 0 diode
R40233 N40232 N40233 10
D40233 N40233 0 diode
R40234 N40233 N40234 10
D40234 N40234 0 diode
R40235 N40234 N40235 10
D40235 N40235 0 diode
R40236 N40235 N40236 10
D40236 N40236 0 diode
R40237 N40236 N40237 10
D40237 N40237 0 diode
R40238 N40237 N40238 10
D40238 N40238 0 diode
R40239 N40238 N40239 10
D40239 N40239 0 diode
R40240 N40239 N40240 10
D40240 N40240 0 diode
R40241 N40240 N40241 10
D40241 N40241 0 diode
R40242 N40241 N40242 10
D40242 N40242 0 diode
R40243 N40242 N40243 10
D40243 N40243 0 diode
R40244 N40243 N40244 10
D40244 N40244 0 diode
R40245 N40244 N40245 10
D40245 N40245 0 diode
R40246 N40245 N40246 10
D40246 N40246 0 diode
R40247 N40246 N40247 10
D40247 N40247 0 diode
R40248 N40247 N40248 10
D40248 N40248 0 diode
R40249 N40248 N40249 10
D40249 N40249 0 diode
R40250 N40249 N40250 10
D40250 N40250 0 diode
R40251 N40250 N40251 10
D40251 N40251 0 diode
R40252 N40251 N40252 10
D40252 N40252 0 diode
R40253 N40252 N40253 10
D40253 N40253 0 diode
R40254 N40253 N40254 10
D40254 N40254 0 diode
R40255 N40254 N40255 10
D40255 N40255 0 diode
R40256 N40255 N40256 10
D40256 N40256 0 diode
R40257 N40256 N40257 10
D40257 N40257 0 diode
R40258 N40257 N40258 10
D40258 N40258 0 diode
R40259 N40258 N40259 10
D40259 N40259 0 diode
R40260 N40259 N40260 10
D40260 N40260 0 diode
R40261 N40260 N40261 10
D40261 N40261 0 diode
R40262 N40261 N40262 10
D40262 N40262 0 diode
R40263 N40262 N40263 10
D40263 N40263 0 diode
R40264 N40263 N40264 10
D40264 N40264 0 diode
R40265 N40264 N40265 10
D40265 N40265 0 diode
R40266 N40265 N40266 10
D40266 N40266 0 diode
R40267 N40266 N40267 10
D40267 N40267 0 diode
R40268 N40267 N40268 10
D40268 N40268 0 diode
R40269 N40268 N40269 10
D40269 N40269 0 diode
R40270 N40269 N40270 10
D40270 N40270 0 diode
R40271 N40270 N40271 10
D40271 N40271 0 diode
R40272 N40271 N40272 10
D40272 N40272 0 diode
R40273 N40272 N40273 10
D40273 N40273 0 diode
R40274 N40273 N40274 10
D40274 N40274 0 diode
R40275 N40274 N40275 10
D40275 N40275 0 diode
R40276 N40275 N40276 10
D40276 N40276 0 diode
R40277 N40276 N40277 10
D40277 N40277 0 diode
R40278 N40277 N40278 10
D40278 N40278 0 diode
R40279 N40278 N40279 10
D40279 N40279 0 diode
R40280 N40279 N40280 10
D40280 N40280 0 diode
R40281 N40280 N40281 10
D40281 N40281 0 diode
R40282 N40281 N40282 10
D40282 N40282 0 diode
R40283 N40282 N40283 10
D40283 N40283 0 diode
R40284 N40283 N40284 10
D40284 N40284 0 diode
R40285 N40284 N40285 10
D40285 N40285 0 diode
R40286 N40285 N40286 10
D40286 N40286 0 diode
R40287 N40286 N40287 10
D40287 N40287 0 diode
R40288 N40287 N40288 10
D40288 N40288 0 diode
R40289 N40288 N40289 10
D40289 N40289 0 diode
R40290 N40289 N40290 10
D40290 N40290 0 diode
R40291 N40290 N40291 10
D40291 N40291 0 diode
R40292 N40291 N40292 10
D40292 N40292 0 diode
R40293 N40292 N40293 10
D40293 N40293 0 diode
R40294 N40293 N40294 10
D40294 N40294 0 diode
R40295 N40294 N40295 10
D40295 N40295 0 diode
R40296 N40295 N40296 10
D40296 N40296 0 diode
R40297 N40296 N40297 10
D40297 N40297 0 diode
R40298 N40297 N40298 10
D40298 N40298 0 diode
R40299 N40298 N40299 10
D40299 N40299 0 diode
R40300 N40299 N40300 10
D40300 N40300 0 diode
R40301 N40300 N40301 10
D40301 N40301 0 diode
R40302 N40301 N40302 10
D40302 N40302 0 diode
R40303 N40302 N40303 10
D40303 N40303 0 diode
R40304 N40303 N40304 10
D40304 N40304 0 diode
R40305 N40304 N40305 10
D40305 N40305 0 diode
R40306 N40305 N40306 10
D40306 N40306 0 diode
R40307 N40306 N40307 10
D40307 N40307 0 diode
R40308 N40307 N40308 10
D40308 N40308 0 diode
R40309 N40308 N40309 10
D40309 N40309 0 diode
R40310 N40309 N40310 10
D40310 N40310 0 diode
R40311 N40310 N40311 10
D40311 N40311 0 diode
R40312 N40311 N40312 10
D40312 N40312 0 diode
R40313 N40312 N40313 10
D40313 N40313 0 diode
R40314 N40313 N40314 10
D40314 N40314 0 diode
R40315 N40314 N40315 10
D40315 N40315 0 diode
R40316 N40315 N40316 10
D40316 N40316 0 diode
R40317 N40316 N40317 10
D40317 N40317 0 diode
R40318 N40317 N40318 10
D40318 N40318 0 diode
R40319 N40318 N40319 10
D40319 N40319 0 diode
R40320 N40319 N40320 10
D40320 N40320 0 diode
R40321 N40320 N40321 10
D40321 N40321 0 diode
R40322 N40321 N40322 10
D40322 N40322 0 diode
R40323 N40322 N40323 10
D40323 N40323 0 diode
R40324 N40323 N40324 10
D40324 N40324 0 diode
R40325 N40324 N40325 10
D40325 N40325 0 diode
R40326 N40325 N40326 10
D40326 N40326 0 diode
R40327 N40326 N40327 10
D40327 N40327 0 diode
R40328 N40327 N40328 10
D40328 N40328 0 diode
R40329 N40328 N40329 10
D40329 N40329 0 diode
R40330 N40329 N40330 10
D40330 N40330 0 diode
R40331 N40330 N40331 10
D40331 N40331 0 diode
R40332 N40331 N40332 10
D40332 N40332 0 diode
R40333 N40332 N40333 10
D40333 N40333 0 diode
R40334 N40333 N40334 10
D40334 N40334 0 diode
R40335 N40334 N40335 10
D40335 N40335 0 diode
R40336 N40335 N40336 10
D40336 N40336 0 diode
R40337 N40336 N40337 10
D40337 N40337 0 diode
R40338 N40337 N40338 10
D40338 N40338 0 diode
R40339 N40338 N40339 10
D40339 N40339 0 diode
R40340 N40339 N40340 10
D40340 N40340 0 diode
R40341 N40340 N40341 10
D40341 N40341 0 diode
R40342 N40341 N40342 10
D40342 N40342 0 diode
R40343 N40342 N40343 10
D40343 N40343 0 diode
R40344 N40343 N40344 10
D40344 N40344 0 diode
R40345 N40344 N40345 10
D40345 N40345 0 diode
R40346 N40345 N40346 10
D40346 N40346 0 diode
R40347 N40346 N40347 10
D40347 N40347 0 diode
R40348 N40347 N40348 10
D40348 N40348 0 diode
R40349 N40348 N40349 10
D40349 N40349 0 diode
R40350 N40349 N40350 10
D40350 N40350 0 diode
R40351 N40350 N40351 10
D40351 N40351 0 diode
R40352 N40351 N40352 10
D40352 N40352 0 diode
R40353 N40352 N40353 10
D40353 N40353 0 diode
R40354 N40353 N40354 10
D40354 N40354 0 diode
R40355 N40354 N40355 10
D40355 N40355 0 diode
R40356 N40355 N40356 10
D40356 N40356 0 diode
R40357 N40356 N40357 10
D40357 N40357 0 diode
R40358 N40357 N40358 10
D40358 N40358 0 diode
R40359 N40358 N40359 10
D40359 N40359 0 diode
R40360 N40359 N40360 10
D40360 N40360 0 diode
R40361 N40360 N40361 10
D40361 N40361 0 diode
R40362 N40361 N40362 10
D40362 N40362 0 diode
R40363 N40362 N40363 10
D40363 N40363 0 diode
R40364 N40363 N40364 10
D40364 N40364 0 diode
R40365 N40364 N40365 10
D40365 N40365 0 diode
R40366 N40365 N40366 10
D40366 N40366 0 diode
R40367 N40366 N40367 10
D40367 N40367 0 diode
R40368 N40367 N40368 10
D40368 N40368 0 diode
R40369 N40368 N40369 10
D40369 N40369 0 diode
R40370 N40369 N40370 10
D40370 N40370 0 diode
R40371 N40370 N40371 10
D40371 N40371 0 diode
R40372 N40371 N40372 10
D40372 N40372 0 diode
R40373 N40372 N40373 10
D40373 N40373 0 diode
R40374 N40373 N40374 10
D40374 N40374 0 diode
R40375 N40374 N40375 10
D40375 N40375 0 diode
R40376 N40375 N40376 10
D40376 N40376 0 diode
R40377 N40376 N40377 10
D40377 N40377 0 diode
R40378 N40377 N40378 10
D40378 N40378 0 diode
R40379 N40378 N40379 10
D40379 N40379 0 diode
R40380 N40379 N40380 10
D40380 N40380 0 diode
R40381 N40380 N40381 10
D40381 N40381 0 diode
R40382 N40381 N40382 10
D40382 N40382 0 diode
R40383 N40382 N40383 10
D40383 N40383 0 diode
R40384 N40383 N40384 10
D40384 N40384 0 diode
R40385 N40384 N40385 10
D40385 N40385 0 diode
R40386 N40385 N40386 10
D40386 N40386 0 diode
R40387 N40386 N40387 10
D40387 N40387 0 diode
R40388 N40387 N40388 10
D40388 N40388 0 diode
R40389 N40388 N40389 10
D40389 N40389 0 diode
R40390 N40389 N40390 10
D40390 N40390 0 diode
R40391 N40390 N40391 10
D40391 N40391 0 diode
R40392 N40391 N40392 10
D40392 N40392 0 diode
R40393 N40392 N40393 10
D40393 N40393 0 diode
R40394 N40393 N40394 10
D40394 N40394 0 diode
R40395 N40394 N40395 10
D40395 N40395 0 diode
R40396 N40395 N40396 10
D40396 N40396 0 diode
R40397 N40396 N40397 10
D40397 N40397 0 diode
R40398 N40397 N40398 10
D40398 N40398 0 diode
R40399 N40398 N40399 10
D40399 N40399 0 diode
R40400 N40399 N40400 10
D40400 N40400 0 diode
R40401 N40400 N40401 10
D40401 N40401 0 diode
R40402 N40401 N40402 10
D40402 N40402 0 diode
R40403 N40402 N40403 10
D40403 N40403 0 diode
R40404 N40403 N40404 10
D40404 N40404 0 diode
R40405 N40404 N40405 10
D40405 N40405 0 diode
R40406 N40405 N40406 10
D40406 N40406 0 diode
R40407 N40406 N40407 10
D40407 N40407 0 diode
R40408 N40407 N40408 10
D40408 N40408 0 diode
R40409 N40408 N40409 10
D40409 N40409 0 diode
R40410 N40409 N40410 10
D40410 N40410 0 diode
R40411 N40410 N40411 10
D40411 N40411 0 diode
R40412 N40411 N40412 10
D40412 N40412 0 diode
R40413 N40412 N40413 10
D40413 N40413 0 diode
R40414 N40413 N40414 10
D40414 N40414 0 diode
R40415 N40414 N40415 10
D40415 N40415 0 diode
R40416 N40415 N40416 10
D40416 N40416 0 diode
R40417 N40416 N40417 10
D40417 N40417 0 diode
R40418 N40417 N40418 10
D40418 N40418 0 diode
R40419 N40418 N40419 10
D40419 N40419 0 diode
R40420 N40419 N40420 10
D40420 N40420 0 diode
R40421 N40420 N40421 10
D40421 N40421 0 diode
R40422 N40421 N40422 10
D40422 N40422 0 diode
R40423 N40422 N40423 10
D40423 N40423 0 diode
R40424 N40423 N40424 10
D40424 N40424 0 diode
R40425 N40424 N40425 10
D40425 N40425 0 diode
R40426 N40425 N40426 10
D40426 N40426 0 diode
R40427 N40426 N40427 10
D40427 N40427 0 diode
R40428 N40427 N40428 10
D40428 N40428 0 diode
R40429 N40428 N40429 10
D40429 N40429 0 diode
R40430 N40429 N40430 10
D40430 N40430 0 diode
R40431 N40430 N40431 10
D40431 N40431 0 diode
R40432 N40431 N40432 10
D40432 N40432 0 diode
R40433 N40432 N40433 10
D40433 N40433 0 diode
R40434 N40433 N40434 10
D40434 N40434 0 diode
R40435 N40434 N40435 10
D40435 N40435 0 diode
R40436 N40435 N40436 10
D40436 N40436 0 diode
R40437 N40436 N40437 10
D40437 N40437 0 diode
R40438 N40437 N40438 10
D40438 N40438 0 diode
R40439 N40438 N40439 10
D40439 N40439 0 diode
R40440 N40439 N40440 10
D40440 N40440 0 diode
R40441 N40440 N40441 10
D40441 N40441 0 diode
R40442 N40441 N40442 10
D40442 N40442 0 diode
R40443 N40442 N40443 10
D40443 N40443 0 diode
R40444 N40443 N40444 10
D40444 N40444 0 diode
R40445 N40444 N40445 10
D40445 N40445 0 diode
R40446 N40445 N40446 10
D40446 N40446 0 diode
R40447 N40446 N40447 10
D40447 N40447 0 diode
R40448 N40447 N40448 10
D40448 N40448 0 diode
R40449 N40448 N40449 10
D40449 N40449 0 diode
R40450 N40449 N40450 10
D40450 N40450 0 diode
R40451 N40450 N40451 10
D40451 N40451 0 diode
R40452 N40451 N40452 10
D40452 N40452 0 diode
R40453 N40452 N40453 10
D40453 N40453 0 diode
R40454 N40453 N40454 10
D40454 N40454 0 diode
R40455 N40454 N40455 10
D40455 N40455 0 diode
R40456 N40455 N40456 10
D40456 N40456 0 diode
R40457 N40456 N40457 10
D40457 N40457 0 diode
R40458 N40457 N40458 10
D40458 N40458 0 diode
R40459 N40458 N40459 10
D40459 N40459 0 diode
R40460 N40459 N40460 10
D40460 N40460 0 diode
R40461 N40460 N40461 10
D40461 N40461 0 diode
R40462 N40461 N40462 10
D40462 N40462 0 diode
R40463 N40462 N40463 10
D40463 N40463 0 diode
R40464 N40463 N40464 10
D40464 N40464 0 diode
R40465 N40464 N40465 10
D40465 N40465 0 diode
R40466 N40465 N40466 10
D40466 N40466 0 diode
R40467 N40466 N40467 10
D40467 N40467 0 diode
R40468 N40467 N40468 10
D40468 N40468 0 diode
R40469 N40468 N40469 10
D40469 N40469 0 diode
R40470 N40469 N40470 10
D40470 N40470 0 diode
R40471 N40470 N40471 10
D40471 N40471 0 diode
R40472 N40471 N40472 10
D40472 N40472 0 diode
R40473 N40472 N40473 10
D40473 N40473 0 diode
R40474 N40473 N40474 10
D40474 N40474 0 diode
R40475 N40474 N40475 10
D40475 N40475 0 diode
R40476 N40475 N40476 10
D40476 N40476 0 diode
R40477 N40476 N40477 10
D40477 N40477 0 diode
R40478 N40477 N40478 10
D40478 N40478 0 diode
R40479 N40478 N40479 10
D40479 N40479 0 diode
R40480 N40479 N40480 10
D40480 N40480 0 diode
R40481 N40480 N40481 10
D40481 N40481 0 diode
R40482 N40481 N40482 10
D40482 N40482 0 diode
R40483 N40482 N40483 10
D40483 N40483 0 diode
R40484 N40483 N40484 10
D40484 N40484 0 diode
R40485 N40484 N40485 10
D40485 N40485 0 diode
R40486 N40485 N40486 10
D40486 N40486 0 diode
R40487 N40486 N40487 10
D40487 N40487 0 diode
R40488 N40487 N40488 10
D40488 N40488 0 diode
R40489 N40488 N40489 10
D40489 N40489 0 diode
R40490 N40489 N40490 10
D40490 N40490 0 diode
R40491 N40490 N40491 10
D40491 N40491 0 diode
R40492 N40491 N40492 10
D40492 N40492 0 diode
R40493 N40492 N40493 10
D40493 N40493 0 diode
R40494 N40493 N40494 10
D40494 N40494 0 diode
R40495 N40494 N40495 10
D40495 N40495 0 diode
R40496 N40495 N40496 10
D40496 N40496 0 diode
R40497 N40496 N40497 10
D40497 N40497 0 diode
R40498 N40497 N40498 10
D40498 N40498 0 diode
R40499 N40498 N40499 10
D40499 N40499 0 diode
R40500 N40499 N40500 10
D40500 N40500 0 diode
R40501 N40500 N40501 10
D40501 N40501 0 diode
R40502 N40501 N40502 10
D40502 N40502 0 diode
R40503 N40502 N40503 10
D40503 N40503 0 diode
R40504 N40503 N40504 10
D40504 N40504 0 diode
R40505 N40504 N40505 10
D40505 N40505 0 diode
R40506 N40505 N40506 10
D40506 N40506 0 diode
R40507 N40506 N40507 10
D40507 N40507 0 diode
R40508 N40507 N40508 10
D40508 N40508 0 diode
R40509 N40508 N40509 10
D40509 N40509 0 diode
R40510 N40509 N40510 10
D40510 N40510 0 diode
R40511 N40510 N40511 10
D40511 N40511 0 diode
R40512 N40511 N40512 10
D40512 N40512 0 diode
R40513 N40512 N40513 10
D40513 N40513 0 diode
R40514 N40513 N40514 10
D40514 N40514 0 diode
R40515 N40514 N40515 10
D40515 N40515 0 diode
R40516 N40515 N40516 10
D40516 N40516 0 diode
R40517 N40516 N40517 10
D40517 N40517 0 diode
R40518 N40517 N40518 10
D40518 N40518 0 diode
R40519 N40518 N40519 10
D40519 N40519 0 diode
R40520 N40519 N40520 10
D40520 N40520 0 diode
R40521 N40520 N40521 10
D40521 N40521 0 diode
R40522 N40521 N40522 10
D40522 N40522 0 diode
R40523 N40522 N40523 10
D40523 N40523 0 diode
R40524 N40523 N40524 10
D40524 N40524 0 diode
R40525 N40524 N40525 10
D40525 N40525 0 diode
R40526 N40525 N40526 10
D40526 N40526 0 diode
R40527 N40526 N40527 10
D40527 N40527 0 diode
R40528 N40527 N40528 10
D40528 N40528 0 diode
R40529 N40528 N40529 10
D40529 N40529 0 diode
R40530 N40529 N40530 10
D40530 N40530 0 diode
R40531 N40530 N40531 10
D40531 N40531 0 diode
R40532 N40531 N40532 10
D40532 N40532 0 diode
R40533 N40532 N40533 10
D40533 N40533 0 diode
R40534 N40533 N40534 10
D40534 N40534 0 diode
R40535 N40534 N40535 10
D40535 N40535 0 diode
R40536 N40535 N40536 10
D40536 N40536 0 diode
R40537 N40536 N40537 10
D40537 N40537 0 diode
R40538 N40537 N40538 10
D40538 N40538 0 diode
R40539 N40538 N40539 10
D40539 N40539 0 diode
R40540 N40539 N40540 10
D40540 N40540 0 diode
R40541 N40540 N40541 10
D40541 N40541 0 diode
R40542 N40541 N40542 10
D40542 N40542 0 diode
R40543 N40542 N40543 10
D40543 N40543 0 diode
R40544 N40543 N40544 10
D40544 N40544 0 diode
R40545 N40544 N40545 10
D40545 N40545 0 diode
R40546 N40545 N40546 10
D40546 N40546 0 diode
R40547 N40546 N40547 10
D40547 N40547 0 diode
R40548 N40547 N40548 10
D40548 N40548 0 diode
R40549 N40548 N40549 10
D40549 N40549 0 diode
R40550 N40549 N40550 10
D40550 N40550 0 diode
R40551 N40550 N40551 10
D40551 N40551 0 diode
R40552 N40551 N40552 10
D40552 N40552 0 diode
R40553 N40552 N40553 10
D40553 N40553 0 diode
R40554 N40553 N40554 10
D40554 N40554 0 diode
R40555 N40554 N40555 10
D40555 N40555 0 diode
R40556 N40555 N40556 10
D40556 N40556 0 diode
R40557 N40556 N40557 10
D40557 N40557 0 diode
R40558 N40557 N40558 10
D40558 N40558 0 diode
R40559 N40558 N40559 10
D40559 N40559 0 diode
R40560 N40559 N40560 10
D40560 N40560 0 diode
R40561 N40560 N40561 10
D40561 N40561 0 diode
R40562 N40561 N40562 10
D40562 N40562 0 diode
R40563 N40562 N40563 10
D40563 N40563 0 diode
R40564 N40563 N40564 10
D40564 N40564 0 diode
R40565 N40564 N40565 10
D40565 N40565 0 diode
R40566 N40565 N40566 10
D40566 N40566 0 diode
R40567 N40566 N40567 10
D40567 N40567 0 diode
R40568 N40567 N40568 10
D40568 N40568 0 diode
R40569 N40568 N40569 10
D40569 N40569 0 diode
R40570 N40569 N40570 10
D40570 N40570 0 diode
R40571 N40570 N40571 10
D40571 N40571 0 diode
R40572 N40571 N40572 10
D40572 N40572 0 diode
R40573 N40572 N40573 10
D40573 N40573 0 diode
R40574 N40573 N40574 10
D40574 N40574 0 diode
R40575 N40574 N40575 10
D40575 N40575 0 diode
R40576 N40575 N40576 10
D40576 N40576 0 diode
R40577 N40576 N40577 10
D40577 N40577 0 diode
R40578 N40577 N40578 10
D40578 N40578 0 diode
R40579 N40578 N40579 10
D40579 N40579 0 diode
R40580 N40579 N40580 10
D40580 N40580 0 diode
R40581 N40580 N40581 10
D40581 N40581 0 diode
R40582 N40581 N40582 10
D40582 N40582 0 diode
R40583 N40582 N40583 10
D40583 N40583 0 diode
R40584 N40583 N40584 10
D40584 N40584 0 diode
R40585 N40584 N40585 10
D40585 N40585 0 diode
R40586 N40585 N40586 10
D40586 N40586 0 diode
R40587 N40586 N40587 10
D40587 N40587 0 diode
R40588 N40587 N40588 10
D40588 N40588 0 diode
R40589 N40588 N40589 10
D40589 N40589 0 diode
R40590 N40589 N40590 10
D40590 N40590 0 diode
R40591 N40590 N40591 10
D40591 N40591 0 diode
R40592 N40591 N40592 10
D40592 N40592 0 diode
R40593 N40592 N40593 10
D40593 N40593 0 diode
R40594 N40593 N40594 10
D40594 N40594 0 diode
R40595 N40594 N40595 10
D40595 N40595 0 diode
R40596 N40595 N40596 10
D40596 N40596 0 diode
R40597 N40596 N40597 10
D40597 N40597 0 diode
R40598 N40597 N40598 10
D40598 N40598 0 diode
R40599 N40598 N40599 10
D40599 N40599 0 diode
R40600 N40599 N40600 10
D40600 N40600 0 diode
R40601 N40600 N40601 10
D40601 N40601 0 diode
R40602 N40601 N40602 10
D40602 N40602 0 diode
R40603 N40602 N40603 10
D40603 N40603 0 diode
R40604 N40603 N40604 10
D40604 N40604 0 diode
R40605 N40604 N40605 10
D40605 N40605 0 diode
R40606 N40605 N40606 10
D40606 N40606 0 diode
R40607 N40606 N40607 10
D40607 N40607 0 diode
R40608 N40607 N40608 10
D40608 N40608 0 diode
R40609 N40608 N40609 10
D40609 N40609 0 diode
R40610 N40609 N40610 10
D40610 N40610 0 diode
R40611 N40610 N40611 10
D40611 N40611 0 diode
R40612 N40611 N40612 10
D40612 N40612 0 diode
R40613 N40612 N40613 10
D40613 N40613 0 diode
R40614 N40613 N40614 10
D40614 N40614 0 diode
R40615 N40614 N40615 10
D40615 N40615 0 diode
R40616 N40615 N40616 10
D40616 N40616 0 diode
R40617 N40616 N40617 10
D40617 N40617 0 diode
R40618 N40617 N40618 10
D40618 N40618 0 diode
R40619 N40618 N40619 10
D40619 N40619 0 diode
R40620 N40619 N40620 10
D40620 N40620 0 diode
R40621 N40620 N40621 10
D40621 N40621 0 diode
R40622 N40621 N40622 10
D40622 N40622 0 diode
R40623 N40622 N40623 10
D40623 N40623 0 diode
R40624 N40623 N40624 10
D40624 N40624 0 diode
R40625 N40624 N40625 10
D40625 N40625 0 diode
R40626 N40625 N40626 10
D40626 N40626 0 diode
R40627 N40626 N40627 10
D40627 N40627 0 diode
R40628 N40627 N40628 10
D40628 N40628 0 diode
R40629 N40628 N40629 10
D40629 N40629 0 diode
R40630 N40629 N40630 10
D40630 N40630 0 diode
R40631 N40630 N40631 10
D40631 N40631 0 diode
R40632 N40631 N40632 10
D40632 N40632 0 diode
R40633 N40632 N40633 10
D40633 N40633 0 diode
R40634 N40633 N40634 10
D40634 N40634 0 diode
R40635 N40634 N40635 10
D40635 N40635 0 diode
R40636 N40635 N40636 10
D40636 N40636 0 diode
R40637 N40636 N40637 10
D40637 N40637 0 diode
R40638 N40637 N40638 10
D40638 N40638 0 diode
R40639 N40638 N40639 10
D40639 N40639 0 diode
R40640 N40639 N40640 10
D40640 N40640 0 diode
R40641 N40640 N40641 10
D40641 N40641 0 diode
R40642 N40641 N40642 10
D40642 N40642 0 diode
R40643 N40642 N40643 10
D40643 N40643 0 diode
R40644 N40643 N40644 10
D40644 N40644 0 diode
R40645 N40644 N40645 10
D40645 N40645 0 diode
R40646 N40645 N40646 10
D40646 N40646 0 diode
R40647 N40646 N40647 10
D40647 N40647 0 diode
R40648 N40647 N40648 10
D40648 N40648 0 diode
R40649 N40648 N40649 10
D40649 N40649 0 diode
R40650 N40649 N40650 10
D40650 N40650 0 diode
R40651 N40650 N40651 10
D40651 N40651 0 diode
R40652 N40651 N40652 10
D40652 N40652 0 diode
R40653 N40652 N40653 10
D40653 N40653 0 diode
R40654 N40653 N40654 10
D40654 N40654 0 diode
R40655 N40654 N40655 10
D40655 N40655 0 diode
R40656 N40655 N40656 10
D40656 N40656 0 diode
R40657 N40656 N40657 10
D40657 N40657 0 diode
R40658 N40657 N40658 10
D40658 N40658 0 diode
R40659 N40658 N40659 10
D40659 N40659 0 diode
R40660 N40659 N40660 10
D40660 N40660 0 diode
R40661 N40660 N40661 10
D40661 N40661 0 diode
R40662 N40661 N40662 10
D40662 N40662 0 diode
R40663 N40662 N40663 10
D40663 N40663 0 diode
R40664 N40663 N40664 10
D40664 N40664 0 diode
R40665 N40664 N40665 10
D40665 N40665 0 diode
R40666 N40665 N40666 10
D40666 N40666 0 diode
R40667 N40666 N40667 10
D40667 N40667 0 diode
R40668 N40667 N40668 10
D40668 N40668 0 diode
R40669 N40668 N40669 10
D40669 N40669 0 diode
R40670 N40669 N40670 10
D40670 N40670 0 diode
R40671 N40670 N40671 10
D40671 N40671 0 diode
R40672 N40671 N40672 10
D40672 N40672 0 diode
R40673 N40672 N40673 10
D40673 N40673 0 diode
R40674 N40673 N40674 10
D40674 N40674 0 diode
R40675 N40674 N40675 10
D40675 N40675 0 diode
R40676 N40675 N40676 10
D40676 N40676 0 diode
R40677 N40676 N40677 10
D40677 N40677 0 diode
R40678 N40677 N40678 10
D40678 N40678 0 diode
R40679 N40678 N40679 10
D40679 N40679 0 diode
R40680 N40679 N40680 10
D40680 N40680 0 diode
R40681 N40680 N40681 10
D40681 N40681 0 diode
R40682 N40681 N40682 10
D40682 N40682 0 diode
R40683 N40682 N40683 10
D40683 N40683 0 diode
R40684 N40683 N40684 10
D40684 N40684 0 diode
R40685 N40684 N40685 10
D40685 N40685 0 diode
R40686 N40685 N40686 10
D40686 N40686 0 diode
R40687 N40686 N40687 10
D40687 N40687 0 diode
R40688 N40687 N40688 10
D40688 N40688 0 diode
R40689 N40688 N40689 10
D40689 N40689 0 diode
R40690 N40689 N40690 10
D40690 N40690 0 diode
R40691 N40690 N40691 10
D40691 N40691 0 diode
R40692 N40691 N40692 10
D40692 N40692 0 diode
R40693 N40692 N40693 10
D40693 N40693 0 diode
R40694 N40693 N40694 10
D40694 N40694 0 diode
R40695 N40694 N40695 10
D40695 N40695 0 diode
R40696 N40695 N40696 10
D40696 N40696 0 diode
R40697 N40696 N40697 10
D40697 N40697 0 diode
R40698 N40697 N40698 10
D40698 N40698 0 diode
R40699 N40698 N40699 10
D40699 N40699 0 diode
R40700 N40699 N40700 10
D40700 N40700 0 diode
R40701 N40700 N40701 10
D40701 N40701 0 diode
R40702 N40701 N40702 10
D40702 N40702 0 diode
R40703 N40702 N40703 10
D40703 N40703 0 diode
R40704 N40703 N40704 10
D40704 N40704 0 diode
R40705 N40704 N40705 10
D40705 N40705 0 diode
R40706 N40705 N40706 10
D40706 N40706 0 diode
R40707 N40706 N40707 10
D40707 N40707 0 diode
R40708 N40707 N40708 10
D40708 N40708 0 diode
R40709 N40708 N40709 10
D40709 N40709 0 diode
R40710 N40709 N40710 10
D40710 N40710 0 diode
R40711 N40710 N40711 10
D40711 N40711 0 diode
R40712 N40711 N40712 10
D40712 N40712 0 diode
R40713 N40712 N40713 10
D40713 N40713 0 diode
R40714 N40713 N40714 10
D40714 N40714 0 diode
R40715 N40714 N40715 10
D40715 N40715 0 diode
R40716 N40715 N40716 10
D40716 N40716 0 diode
R40717 N40716 N40717 10
D40717 N40717 0 diode
R40718 N40717 N40718 10
D40718 N40718 0 diode
R40719 N40718 N40719 10
D40719 N40719 0 diode
R40720 N40719 N40720 10
D40720 N40720 0 diode
R40721 N40720 N40721 10
D40721 N40721 0 diode
R40722 N40721 N40722 10
D40722 N40722 0 diode
R40723 N40722 N40723 10
D40723 N40723 0 diode
R40724 N40723 N40724 10
D40724 N40724 0 diode
R40725 N40724 N40725 10
D40725 N40725 0 diode
R40726 N40725 N40726 10
D40726 N40726 0 diode
R40727 N40726 N40727 10
D40727 N40727 0 diode
R40728 N40727 N40728 10
D40728 N40728 0 diode
R40729 N40728 N40729 10
D40729 N40729 0 diode
R40730 N40729 N40730 10
D40730 N40730 0 diode
R40731 N40730 N40731 10
D40731 N40731 0 diode
R40732 N40731 N40732 10
D40732 N40732 0 diode
R40733 N40732 N40733 10
D40733 N40733 0 diode
R40734 N40733 N40734 10
D40734 N40734 0 diode
R40735 N40734 N40735 10
D40735 N40735 0 diode
R40736 N40735 N40736 10
D40736 N40736 0 diode
R40737 N40736 N40737 10
D40737 N40737 0 diode
R40738 N40737 N40738 10
D40738 N40738 0 diode
R40739 N40738 N40739 10
D40739 N40739 0 diode
R40740 N40739 N40740 10
D40740 N40740 0 diode
R40741 N40740 N40741 10
D40741 N40741 0 diode
R40742 N40741 N40742 10
D40742 N40742 0 diode
R40743 N40742 N40743 10
D40743 N40743 0 diode
R40744 N40743 N40744 10
D40744 N40744 0 diode
R40745 N40744 N40745 10
D40745 N40745 0 diode
R40746 N40745 N40746 10
D40746 N40746 0 diode
R40747 N40746 N40747 10
D40747 N40747 0 diode
R40748 N40747 N40748 10
D40748 N40748 0 diode
R40749 N40748 N40749 10
D40749 N40749 0 diode
R40750 N40749 N40750 10
D40750 N40750 0 diode
R40751 N40750 N40751 10
D40751 N40751 0 diode
R40752 N40751 N40752 10
D40752 N40752 0 diode
R40753 N40752 N40753 10
D40753 N40753 0 diode
R40754 N40753 N40754 10
D40754 N40754 0 diode
R40755 N40754 N40755 10
D40755 N40755 0 diode
R40756 N40755 N40756 10
D40756 N40756 0 diode
R40757 N40756 N40757 10
D40757 N40757 0 diode
R40758 N40757 N40758 10
D40758 N40758 0 diode
R40759 N40758 N40759 10
D40759 N40759 0 diode
R40760 N40759 N40760 10
D40760 N40760 0 diode
R40761 N40760 N40761 10
D40761 N40761 0 diode
R40762 N40761 N40762 10
D40762 N40762 0 diode
R40763 N40762 N40763 10
D40763 N40763 0 diode
R40764 N40763 N40764 10
D40764 N40764 0 diode
R40765 N40764 N40765 10
D40765 N40765 0 diode
R40766 N40765 N40766 10
D40766 N40766 0 diode
R40767 N40766 N40767 10
D40767 N40767 0 diode
R40768 N40767 N40768 10
D40768 N40768 0 diode
R40769 N40768 N40769 10
D40769 N40769 0 diode
R40770 N40769 N40770 10
D40770 N40770 0 diode
R40771 N40770 N40771 10
D40771 N40771 0 diode
R40772 N40771 N40772 10
D40772 N40772 0 diode
R40773 N40772 N40773 10
D40773 N40773 0 diode
R40774 N40773 N40774 10
D40774 N40774 0 diode
R40775 N40774 N40775 10
D40775 N40775 0 diode
R40776 N40775 N40776 10
D40776 N40776 0 diode
R40777 N40776 N40777 10
D40777 N40777 0 diode
R40778 N40777 N40778 10
D40778 N40778 0 diode
R40779 N40778 N40779 10
D40779 N40779 0 diode
R40780 N40779 N40780 10
D40780 N40780 0 diode
R40781 N40780 N40781 10
D40781 N40781 0 diode
R40782 N40781 N40782 10
D40782 N40782 0 diode
R40783 N40782 N40783 10
D40783 N40783 0 diode
R40784 N40783 N40784 10
D40784 N40784 0 diode
R40785 N40784 N40785 10
D40785 N40785 0 diode
R40786 N40785 N40786 10
D40786 N40786 0 diode
R40787 N40786 N40787 10
D40787 N40787 0 diode
R40788 N40787 N40788 10
D40788 N40788 0 diode
R40789 N40788 N40789 10
D40789 N40789 0 diode
R40790 N40789 N40790 10
D40790 N40790 0 diode
R40791 N40790 N40791 10
D40791 N40791 0 diode
R40792 N40791 N40792 10
D40792 N40792 0 diode
R40793 N40792 N40793 10
D40793 N40793 0 diode
R40794 N40793 N40794 10
D40794 N40794 0 diode
R40795 N40794 N40795 10
D40795 N40795 0 diode
R40796 N40795 N40796 10
D40796 N40796 0 diode
R40797 N40796 N40797 10
D40797 N40797 0 diode
R40798 N40797 N40798 10
D40798 N40798 0 diode
R40799 N40798 N40799 10
D40799 N40799 0 diode
R40800 N40799 N40800 10
D40800 N40800 0 diode
R40801 N40800 N40801 10
D40801 N40801 0 diode
R40802 N40801 N40802 10
D40802 N40802 0 diode
R40803 N40802 N40803 10
D40803 N40803 0 diode
R40804 N40803 N40804 10
D40804 N40804 0 diode
R40805 N40804 N40805 10
D40805 N40805 0 diode
R40806 N40805 N40806 10
D40806 N40806 0 diode
R40807 N40806 N40807 10
D40807 N40807 0 diode
R40808 N40807 N40808 10
D40808 N40808 0 diode
R40809 N40808 N40809 10
D40809 N40809 0 diode
R40810 N40809 N40810 10
D40810 N40810 0 diode
R40811 N40810 N40811 10
D40811 N40811 0 diode
R40812 N40811 N40812 10
D40812 N40812 0 diode
R40813 N40812 N40813 10
D40813 N40813 0 diode
R40814 N40813 N40814 10
D40814 N40814 0 diode
R40815 N40814 N40815 10
D40815 N40815 0 diode
R40816 N40815 N40816 10
D40816 N40816 0 diode
R40817 N40816 N40817 10
D40817 N40817 0 diode
R40818 N40817 N40818 10
D40818 N40818 0 diode
R40819 N40818 N40819 10
D40819 N40819 0 diode
R40820 N40819 N40820 10
D40820 N40820 0 diode
R40821 N40820 N40821 10
D40821 N40821 0 diode
R40822 N40821 N40822 10
D40822 N40822 0 diode
R40823 N40822 N40823 10
D40823 N40823 0 diode
R40824 N40823 N40824 10
D40824 N40824 0 diode
R40825 N40824 N40825 10
D40825 N40825 0 diode
R40826 N40825 N40826 10
D40826 N40826 0 diode
R40827 N40826 N40827 10
D40827 N40827 0 diode
R40828 N40827 N40828 10
D40828 N40828 0 diode
R40829 N40828 N40829 10
D40829 N40829 0 diode
R40830 N40829 N40830 10
D40830 N40830 0 diode
R40831 N40830 N40831 10
D40831 N40831 0 diode
R40832 N40831 N40832 10
D40832 N40832 0 diode
R40833 N40832 N40833 10
D40833 N40833 0 diode
R40834 N40833 N40834 10
D40834 N40834 0 diode
R40835 N40834 N40835 10
D40835 N40835 0 diode
R40836 N40835 N40836 10
D40836 N40836 0 diode
R40837 N40836 N40837 10
D40837 N40837 0 diode
R40838 N40837 N40838 10
D40838 N40838 0 diode
R40839 N40838 N40839 10
D40839 N40839 0 diode
R40840 N40839 N40840 10
D40840 N40840 0 diode
R40841 N40840 N40841 10
D40841 N40841 0 diode
R40842 N40841 N40842 10
D40842 N40842 0 diode
R40843 N40842 N40843 10
D40843 N40843 0 diode
R40844 N40843 N40844 10
D40844 N40844 0 diode
R40845 N40844 N40845 10
D40845 N40845 0 diode
R40846 N40845 N40846 10
D40846 N40846 0 diode
R40847 N40846 N40847 10
D40847 N40847 0 diode
R40848 N40847 N40848 10
D40848 N40848 0 diode
R40849 N40848 N40849 10
D40849 N40849 0 diode
R40850 N40849 N40850 10
D40850 N40850 0 diode
R40851 N40850 N40851 10
D40851 N40851 0 diode
R40852 N40851 N40852 10
D40852 N40852 0 diode
R40853 N40852 N40853 10
D40853 N40853 0 diode
R40854 N40853 N40854 10
D40854 N40854 0 diode
R40855 N40854 N40855 10
D40855 N40855 0 diode
R40856 N40855 N40856 10
D40856 N40856 0 diode
R40857 N40856 N40857 10
D40857 N40857 0 diode
R40858 N40857 N40858 10
D40858 N40858 0 diode
R40859 N40858 N40859 10
D40859 N40859 0 diode
R40860 N40859 N40860 10
D40860 N40860 0 diode
R40861 N40860 N40861 10
D40861 N40861 0 diode
R40862 N40861 N40862 10
D40862 N40862 0 diode
R40863 N40862 N40863 10
D40863 N40863 0 diode
R40864 N40863 N40864 10
D40864 N40864 0 diode
R40865 N40864 N40865 10
D40865 N40865 0 diode
R40866 N40865 N40866 10
D40866 N40866 0 diode
R40867 N40866 N40867 10
D40867 N40867 0 diode
R40868 N40867 N40868 10
D40868 N40868 0 diode
R40869 N40868 N40869 10
D40869 N40869 0 diode
R40870 N40869 N40870 10
D40870 N40870 0 diode
R40871 N40870 N40871 10
D40871 N40871 0 diode
R40872 N40871 N40872 10
D40872 N40872 0 diode
R40873 N40872 N40873 10
D40873 N40873 0 diode
R40874 N40873 N40874 10
D40874 N40874 0 diode
R40875 N40874 N40875 10
D40875 N40875 0 diode
R40876 N40875 N40876 10
D40876 N40876 0 diode
R40877 N40876 N40877 10
D40877 N40877 0 diode
R40878 N40877 N40878 10
D40878 N40878 0 diode
R40879 N40878 N40879 10
D40879 N40879 0 diode
R40880 N40879 N40880 10
D40880 N40880 0 diode
R40881 N40880 N40881 10
D40881 N40881 0 diode
R40882 N40881 N40882 10
D40882 N40882 0 diode
R40883 N40882 N40883 10
D40883 N40883 0 diode
R40884 N40883 N40884 10
D40884 N40884 0 diode
R40885 N40884 N40885 10
D40885 N40885 0 diode
R40886 N40885 N40886 10
D40886 N40886 0 diode
R40887 N40886 N40887 10
D40887 N40887 0 diode
R40888 N40887 N40888 10
D40888 N40888 0 diode
R40889 N40888 N40889 10
D40889 N40889 0 diode
R40890 N40889 N40890 10
D40890 N40890 0 diode
R40891 N40890 N40891 10
D40891 N40891 0 diode
R40892 N40891 N40892 10
D40892 N40892 0 diode
R40893 N40892 N40893 10
D40893 N40893 0 diode
R40894 N40893 N40894 10
D40894 N40894 0 diode
R40895 N40894 N40895 10
D40895 N40895 0 diode
R40896 N40895 N40896 10
D40896 N40896 0 diode
R40897 N40896 N40897 10
D40897 N40897 0 diode
R40898 N40897 N40898 10
D40898 N40898 0 diode
R40899 N40898 N40899 10
D40899 N40899 0 diode
R40900 N40899 N40900 10
D40900 N40900 0 diode
R40901 N40900 N40901 10
D40901 N40901 0 diode
R40902 N40901 N40902 10
D40902 N40902 0 diode
R40903 N40902 N40903 10
D40903 N40903 0 diode
R40904 N40903 N40904 10
D40904 N40904 0 diode
R40905 N40904 N40905 10
D40905 N40905 0 diode
R40906 N40905 N40906 10
D40906 N40906 0 diode
R40907 N40906 N40907 10
D40907 N40907 0 diode
R40908 N40907 N40908 10
D40908 N40908 0 diode
R40909 N40908 N40909 10
D40909 N40909 0 diode
R40910 N40909 N40910 10
D40910 N40910 0 diode
R40911 N40910 N40911 10
D40911 N40911 0 diode
R40912 N40911 N40912 10
D40912 N40912 0 diode
R40913 N40912 N40913 10
D40913 N40913 0 diode
R40914 N40913 N40914 10
D40914 N40914 0 diode
R40915 N40914 N40915 10
D40915 N40915 0 diode
R40916 N40915 N40916 10
D40916 N40916 0 diode
R40917 N40916 N40917 10
D40917 N40917 0 diode
R40918 N40917 N40918 10
D40918 N40918 0 diode
R40919 N40918 N40919 10
D40919 N40919 0 diode
R40920 N40919 N40920 10
D40920 N40920 0 diode
R40921 N40920 N40921 10
D40921 N40921 0 diode
R40922 N40921 N40922 10
D40922 N40922 0 diode
R40923 N40922 N40923 10
D40923 N40923 0 diode
R40924 N40923 N40924 10
D40924 N40924 0 diode
R40925 N40924 N40925 10
D40925 N40925 0 diode
R40926 N40925 N40926 10
D40926 N40926 0 diode
R40927 N40926 N40927 10
D40927 N40927 0 diode
R40928 N40927 N40928 10
D40928 N40928 0 diode
R40929 N40928 N40929 10
D40929 N40929 0 diode
R40930 N40929 N40930 10
D40930 N40930 0 diode
R40931 N40930 N40931 10
D40931 N40931 0 diode
R40932 N40931 N40932 10
D40932 N40932 0 diode
R40933 N40932 N40933 10
D40933 N40933 0 diode
R40934 N40933 N40934 10
D40934 N40934 0 diode
R40935 N40934 N40935 10
D40935 N40935 0 diode
R40936 N40935 N40936 10
D40936 N40936 0 diode
R40937 N40936 N40937 10
D40937 N40937 0 diode
R40938 N40937 N40938 10
D40938 N40938 0 diode
R40939 N40938 N40939 10
D40939 N40939 0 diode
R40940 N40939 N40940 10
D40940 N40940 0 diode
R40941 N40940 N40941 10
D40941 N40941 0 diode
R40942 N40941 N40942 10
D40942 N40942 0 diode
R40943 N40942 N40943 10
D40943 N40943 0 diode
R40944 N40943 N40944 10
D40944 N40944 0 diode
R40945 N40944 N40945 10
D40945 N40945 0 diode
R40946 N40945 N40946 10
D40946 N40946 0 diode
R40947 N40946 N40947 10
D40947 N40947 0 diode
R40948 N40947 N40948 10
D40948 N40948 0 diode
R40949 N40948 N40949 10
D40949 N40949 0 diode
R40950 N40949 N40950 10
D40950 N40950 0 diode
R40951 N40950 N40951 10
D40951 N40951 0 diode
R40952 N40951 N40952 10
D40952 N40952 0 diode
R40953 N40952 N40953 10
D40953 N40953 0 diode
R40954 N40953 N40954 10
D40954 N40954 0 diode
R40955 N40954 N40955 10
D40955 N40955 0 diode
R40956 N40955 N40956 10
D40956 N40956 0 diode
R40957 N40956 N40957 10
D40957 N40957 0 diode
R40958 N40957 N40958 10
D40958 N40958 0 diode
R40959 N40958 N40959 10
D40959 N40959 0 diode
R40960 N40959 N40960 10
D40960 N40960 0 diode
R40961 N40960 N40961 10
D40961 N40961 0 diode
R40962 N40961 N40962 10
D40962 N40962 0 diode
R40963 N40962 N40963 10
D40963 N40963 0 diode
R40964 N40963 N40964 10
D40964 N40964 0 diode
R40965 N40964 N40965 10
D40965 N40965 0 diode
R40966 N40965 N40966 10
D40966 N40966 0 diode
R40967 N40966 N40967 10
D40967 N40967 0 diode
R40968 N40967 N40968 10
D40968 N40968 0 diode
R40969 N40968 N40969 10
D40969 N40969 0 diode
R40970 N40969 N40970 10
D40970 N40970 0 diode
R40971 N40970 N40971 10
D40971 N40971 0 diode
R40972 N40971 N40972 10
D40972 N40972 0 diode
R40973 N40972 N40973 10
D40973 N40973 0 diode
R40974 N40973 N40974 10
D40974 N40974 0 diode
R40975 N40974 N40975 10
D40975 N40975 0 diode
R40976 N40975 N40976 10
D40976 N40976 0 diode
R40977 N40976 N40977 10
D40977 N40977 0 diode
R40978 N40977 N40978 10
D40978 N40978 0 diode
R40979 N40978 N40979 10
D40979 N40979 0 diode
R40980 N40979 N40980 10
D40980 N40980 0 diode
R40981 N40980 N40981 10
D40981 N40981 0 diode
R40982 N40981 N40982 10
D40982 N40982 0 diode
R40983 N40982 N40983 10
D40983 N40983 0 diode
R40984 N40983 N40984 10
D40984 N40984 0 diode
R40985 N40984 N40985 10
D40985 N40985 0 diode
R40986 N40985 N40986 10
D40986 N40986 0 diode
R40987 N40986 N40987 10
D40987 N40987 0 diode
R40988 N40987 N40988 10
D40988 N40988 0 diode
R40989 N40988 N40989 10
D40989 N40989 0 diode
R40990 N40989 N40990 10
D40990 N40990 0 diode
R40991 N40990 N40991 10
D40991 N40991 0 diode
R40992 N40991 N40992 10
D40992 N40992 0 diode
R40993 N40992 N40993 10
D40993 N40993 0 diode
R40994 N40993 N40994 10
D40994 N40994 0 diode
R40995 N40994 N40995 10
D40995 N40995 0 diode
R40996 N40995 N40996 10
D40996 N40996 0 diode
R40997 N40996 N40997 10
D40997 N40997 0 diode
R40998 N40997 N40998 10
D40998 N40998 0 diode
R40999 N40998 N40999 10
D40999 N40999 0 diode
R41000 N40999 N41000 10
D41000 N41000 0 diode
R41001 N41000 N41001 10
D41001 N41001 0 diode
R41002 N41001 N41002 10
D41002 N41002 0 diode
R41003 N41002 N41003 10
D41003 N41003 0 diode
R41004 N41003 N41004 10
D41004 N41004 0 diode
R41005 N41004 N41005 10
D41005 N41005 0 diode
R41006 N41005 N41006 10
D41006 N41006 0 diode
R41007 N41006 N41007 10
D41007 N41007 0 diode
R41008 N41007 N41008 10
D41008 N41008 0 diode
R41009 N41008 N41009 10
D41009 N41009 0 diode
R41010 N41009 N41010 10
D41010 N41010 0 diode
R41011 N41010 N41011 10
D41011 N41011 0 diode
R41012 N41011 N41012 10
D41012 N41012 0 diode
R41013 N41012 N41013 10
D41013 N41013 0 diode
R41014 N41013 N41014 10
D41014 N41014 0 diode
R41015 N41014 N41015 10
D41015 N41015 0 diode
R41016 N41015 N41016 10
D41016 N41016 0 diode
R41017 N41016 N41017 10
D41017 N41017 0 diode
R41018 N41017 N41018 10
D41018 N41018 0 diode
R41019 N41018 N41019 10
D41019 N41019 0 diode
R41020 N41019 N41020 10
D41020 N41020 0 diode
R41021 N41020 N41021 10
D41021 N41021 0 diode
R41022 N41021 N41022 10
D41022 N41022 0 diode
R41023 N41022 N41023 10
D41023 N41023 0 diode
R41024 N41023 N41024 10
D41024 N41024 0 diode
R41025 N41024 N41025 10
D41025 N41025 0 diode
R41026 N41025 N41026 10
D41026 N41026 0 diode
R41027 N41026 N41027 10
D41027 N41027 0 diode
R41028 N41027 N41028 10
D41028 N41028 0 diode
R41029 N41028 N41029 10
D41029 N41029 0 diode
R41030 N41029 N41030 10
D41030 N41030 0 diode
R41031 N41030 N41031 10
D41031 N41031 0 diode
R41032 N41031 N41032 10
D41032 N41032 0 diode
R41033 N41032 N41033 10
D41033 N41033 0 diode
R41034 N41033 N41034 10
D41034 N41034 0 diode
R41035 N41034 N41035 10
D41035 N41035 0 diode
R41036 N41035 N41036 10
D41036 N41036 0 diode
R41037 N41036 N41037 10
D41037 N41037 0 diode
R41038 N41037 N41038 10
D41038 N41038 0 diode
R41039 N41038 N41039 10
D41039 N41039 0 diode
R41040 N41039 N41040 10
D41040 N41040 0 diode
R41041 N41040 N41041 10
D41041 N41041 0 diode
R41042 N41041 N41042 10
D41042 N41042 0 diode
R41043 N41042 N41043 10
D41043 N41043 0 diode
R41044 N41043 N41044 10
D41044 N41044 0 diode
R41045 N41044 N41045 10
D41045 N41045 0 diode
R41046 N41045 N41046 10
D41046 N41046 0 diode
R41047 N41046 N41047 10
D41047 N41047 0 diode
R41048 N41047 N41048 10
D41048 N41048 0 diode
R41049 N41048 N41049 10
D41049 N41049 0 diode
R41050 N41049 N41050 10
D41050 N41050 0 diode
R41051 N41050 N41051 10
D41051 N41051 0 diode
R41052 N41051 N41052 10
D41052 N41052 0 diode
R41053 N41052 N41053 10
D41053 N41053 0 diode
R41054 N41053 N41054 10
D41054 N41054 0 diode
R41055 N41054 N41055 10
D41055 N41055 0 diode
R41056 N41055 N41056 10
D41056 N41056 0 diode
R41057 N41056 N41057 10
D41057 N41057 0 diode
R41058 N41057 N41058 10
D41058 N41058 0 diode
R41059 N41058 N41059 10
D41059 N41059 0 diode
R41060 N41059 N41060 10
D41060 N41060 0 diode
R41061 N41060 N41061 10
D41061 N41061 0 diode
R41062 N41061 N41062 10
D41062 N41062 0 diode
R41063 N41062 N41063 10
D41063 N41063 0 diode
R41064 N41063 N41064 10
D41064 N41064 0 diode
R41065 N41064 N41065 10
D41065 N41065 0 diode
R41066 N41065 N41066 10
D41066 N41066 0 diode
R41067 N41066 N41067 10
D41067 N41067 0 diode
R41068 N41067 N41068 10
D41068 N41068 0 diode
R41069 N41068 N41069 10
D41069 N41069 0 diode
R41070 N41069 N41070 10
D41070 N41070 0 diode
R41071 N41070 N41071 10
D41071 N41071 0 diode
R41072 N41071 N41072 10
D41072 N41072 0 diode
R41073 N41072 N41073 10
D41073 N41073 0 diode
R41074 N41073 N41074 10
D41074 N41074 0 diode
R41075 N41074 N41075 10
D41075 N41075 0 diode
R41076 N41075 N41076 10
D41076 N41076 0 diode
R41077 N41076 N41077 10
D41077 N41077 0 diode
R41078 N41077 N41078 10
D41078 N41078 0 diode
R41079 N41078 N41079 10
D41079 N41079 0 diode
R41080 N41079 N41080 10
D41080 N41080 0 diode
R41081 N41080 N41081 10
D41081 N41081 0 diode
R41082 N41081 N41082 10
D41082 N41082 0 diode
R41083 N41082 N41083 10
D41083 N41083 0 diode
R41084 N41083 N41084 10
D41084 N41084 0 diode
R41085 N41084 N41085 10
D41085 N41085 0 diode
R41086 N41085 N41086 10
D41086 N41086 0 diode
R41087 N41086 N41087 10
D41087 N41087 0 diode
R41088 N41087 N41088 10
D41088 N41088 0 diode
R41089 N41088 N41089 10
D41089 N41089 0 diode
R41090 N41089 N41090 10
D41090 N41090 0 diode
R41091 N41090 N41091 10
D41091 N41091 0 diode
R41092 N41091 N41092 10
D41092 N41092 0 diode
R41093 N41092 N41093 10
D41093 N41093 0 diode
R41094 N41093 N41094 10
D41094 N41094 0 diode
R41095 N41094 N41095 10
D41095 N41095 0 diode
R41096 N41095 N41096 10
D41096 N41096 0 diode
R41097 N41096 N41097 10
D41097 N41097 0 diode
R41098 N41097 N41098 10
D41098 N41098 0 diode
R41099 N41098 N41099 10
D41099 N41099 0 diode
R41100 N41099 N41100 10
D41100 N41100 0 diode
R41101 N41100 N41101 10
D41101 N41101 0 diode
R41102 N41101 N41102 10
D41102 N41102 0 diode
R41103 N41102 N41103 10
D41103 N41103 0 diode
R41104 N41103 N41104 10
D41104 N41104 0 diode
R41105 N41104 N41105 10
D41105 N41105 0 diode
R41106 N41105 N41106 10
D41106 N41106 0 diode
R41107 N41106 N41107 10
D41107 N41107 0 diode
R41108 N41107 N41108 10
D41108 N41108 0 diode
R41109 N41108 N41109 10
D41109 N41109 0 diode
R41110 N41109 N41110 10
D41110 N41110 0 diode
R41111 N41110 N41111 10
D41111 N41111 0 diode
R41112 N41111 N41112 10
D41112 N41112 0 diode
R41113 N41112 N41113 10
D41113 N41113 0 diode
R41114 N41113 N41114 10
D41114 N41114 0 diode
R41115 N41114 N41115 10
D41115 N41115 0 diode
R41116 N41115 N41116 10
D41116 N41116 0 diode
R41117 N41116 N41117 10
D41117 N41117 0 diode
R41118 N41117 N41118 10
D41118 N41118 0 diode
R41119 N41118 N41119 10
D41119 N41119 0 diode
R41120 N41119 N41120 10
D41120 N41120 0 diode
R41121 N41120 N41121 10
D41121 N41121 0 diode
R41122 N41121 N41122 10
D41122 N41122 0 diode
R41123 N41122 N41123 10
D41123 N41123 0 diode
R41124 N41123 N41124 10
D41124 N41124 0 diode
R41125 N41124 N41125 10
D41125 N41125 0 diode
R41126 N41125 N41126 10
D41126 N41126 0 diode
R41127 N41126 N41127 10
D41127 N41127 0 diode
R41128 N41127 N41128 10
D41128 N41128 0 diode
R41129 N41128 N41129 10
D41129 N41129 0 diode
R41130 N41129 N41130 10
D41130 N41130 0 diode
R41131 N41130 N41131 10
D41131 N41131 0 diode
R41132 N41131 N41132 10
D41132 N41132 0 diode
R41133 N41132 N41133 10
D41133 N41133 0 diode
R41134 N41133 N41134 10
D41134 N41134 0 diode
R41135 N41134 N41135 10
D41135 N41135 0 diode
R41136 N41135 N41136 10
D41136 N41136 0 diode
R41137 N41136 N41137 10
D41137 N41137 0 diode
R41138 N41137 N41138 10
D41138 N41138 0 diode
R41139 N41138 N41139 10
D41139 N41139 0 diode
R41140 N41139 N41140 10
D41140 N41140 0 diode
R41141 N41140 N41141 10
D41141 N41141 0 diode
R41142 N41141 N41142 10
D41142 N41142 0 diode
R41143 N41142 N41143 10
D41143 N41143 0 diode
R41144 N41143 N41144 10
D41144 N41144 0 diode
R41145 N41144 N41145 10
D41145 N41145 0 diode
R41146 N41145 N41146 10
D41146 N41146 0 diode
R41147 N41146 N41147 10
D41147 N41147 0 diode
R41148 N41147 N41148 10
D41148 N41148 0 diode
R41149 N41148 N41149 10
D41149 N41149 0 diode
R41150 N41149 N41150 10
D41150 N41150 0 diode
R41151 N41150 N41151 10
D41151 N41151 0 diode
R41152 N41151 N41152 10
D41152 N41152 0 diode
R41153 N41152 N41153 10
D41153 N41153 0 diode
R41154 N41153 N41154 10
D41154 N41154 0 diode
R41155 N41154 N41155 10
D41155 N41155 0 diode
R41156 N41155 N41156 10
D41156 N41156 0 diode
R41157 N41156 N41157 10
D41157 N41157 0 diode
R41158 N41157 N41158 10
D41158 N41158 0 diode
R41159 N41158 N41159 10
D41159 N41159 0 diode
R41160 N41159 N41160 10
D41160 N41160 0 diode
R41161 N41160 N41161 10
D41161 N41161 0 diode
R41162 N41161 N41162 10
D41162 N41162 0 diode
R41163 N41162 N41163 10
D41163 N41163 0 diode
R41164 N41163 N41164 10
D41164 N41164 0 diode
R41165 N41164 N41165 10
D41165 N41165 0 diode
R41166 N41165 N41166 10
D41166 N41166 0 diode
R41167 N41166 N41167 10
D41167 N41167 0 diode
R41168 N41167 N41168 10
D41168 N41168 0 diode
R41169 N41168 N41169 10
D41169 N41169 0 diode
R41170 N41169 N41170 10
D41170 N41170 0 diode
R41171 N41170 N41171 10
D41171 N41171 0 diode
R41172 N41171 N41172 10
D41172 N41172 0 diode
R41173 N41172 N41173 10
D41173 N41173 0 diode
R41174 N41173 N41174 10
D41174 N41174 0 diode
R41175 N41174 N41175 10
D41175 N41175 0 diode
R41176 N41175 N41176 10
D41176 N41176 0 diode
R41177 N41176 N41177 10
D41177 N41177 0 diode
R41178 N41177 N41178 10
D41178 N41178 0 diode
R41179 N41178 N41179 10
D41179 N41179 0 diode
R41180 N41179 N41180 10
D41180 N41180 0 diode
R41181 N41180 N41181 10
D41181 N41181 0 diode
R41182 N41181 N41182 10
D41182 N41182 0 diode
R41183 N41182 N41183 10
D41183 N41183 0 diode
R41184 N41183 N41184 10
D41184 N41184 0 diode
R41185 N41184 N41185 10
D41185 N41185 0 diode
R41186 N41185 N41186 10
D41186 N41186 0 diode
R41187 N41186 N41187 10
D41187 N41187 0 diode
R41188 N41187 N41188 10
D41188 N41188 0 diode
R41189 N41188 N41189 10
D41189 N41189 0 diode
R41190 N41189 N41190 10
D41190 N41190 0 diode
R41191 N41190 N41191 10
D41191 N41191 0 diode
R41192 N41191 N41192 10
D41192 N41192 0 diode
R41193 N41192 N41193 10
D41193 N41193 0 diode
R41194 N41193 N41194 10
D41194 N41194 0 diode
R41195 N41194 N41195 10
D41195 N41195 0 diode
R41196 N41195 N41196 10
D41196 N41196 0 diode
R41197 N41196 N41197 10
D41197 N41197 0 diode
R41198 N41197 N41198 10
D41198 N41198 0 diode
R41199 N41198 N41199 10
D41199 N41199 0 diode
R41200 N41199 N41200 10
D41200 N41200 0 diode
R41201 N41200 N41201 10
D41201 N41201 0 diode
R41202 N41201 N41202 10
D41202 N41202 0 diode
R41203 N41202 N41203 10
D41203 N41203 0 diode
R41204 N41203 N41204 10
D41204 N41204 0 diode
R41205 N41204 N41205 10
D41205 N41205 0 diode
R41206 N41205 N41206 10
D41206 N41206 0 diode
R41207 N41206 N41207 10
D41207 N41207 0 diode
R41208 N41207 N41208 10
D41208 N41208 0 diode
R41209 N41208 N41209 10
D41209 N41209 0 diode
R41210 N41209 N41210 10
D41210 N41210 0 diode
R41211 N41210 N41211 10
D41211 N41211 0 diode
R41212 N41211 N41212 10
D41212 N41212 0 diode
R41213 N41212 N41213 10
D41213 N41213 0 diode
R41214 N41213 N41214 10
D41214 N41214 0 diode
R41215 N41214 N41215 10
D41215 N41215 0 diode
R41216 N41215 N41216 10
D41216 N41216 0 diode
R41217 N41216 N41217 10
D41217 N41217 0 diode
R41218 N41217 N41218 10
D41218 N41218 0 diode
R41219 N41218 N41219 10
D41219 N41219 0 diode
R41220 N41219 N41220 10
D41220 N41220 0 diode
R41221 N41220 N41221 10
D41221 N41221 0 diode
R41222 N41221 N41222 10
D41222 N41222 0 diode
R41223 N41222 N41223 10
D41223 N41223 0 diode
R41224 N41223 N41224 10
D41224 N41224 0 diode
R41225 N41224 N41225 10
D41225 N41225 0 diode
R41226 N41225 N41226 10
D41226 N41226 0 diode
R41227 N41226 N41227 10
D41227 N41227 0 diode
R41228 N41227 N41228 10
D41228 N41228 0 diode
R41229 N41228 N41229 10
D41229 N41229 0 diode
R41230 N41229 N41230 10
D41230 N41230 0 diode
R41231 N41230 N41231 10
D41231 N41231 0 diode
R41232 N41231 N41232 10
D41232 N41232 0 diode
R41233 N41232 N41233 10
D41233 N41233 0 diode
R41234 N41233 N41234 10
D41234 N41234 0 diode
R41235 N41234 N41235 10
D41235 N41235 0 diode
R41236 N41235 N41236 10
D41236 N41236 0 diode
R41237 N41236 N41237 10
D41237 N41237 0 diode
R41238 N41237 N41238 10
D41238 N41238 0 diode
R41239 N41238 N41239 10
D41239 N41239 0 diode
R41240 N41239 N41240 10
D41240 N41240 0 diode
R41241 N41240 N41241 10
D41241 N41241 0 diode
R41242 N41241 N41242 10
D41242 N41242 0 diode
R41243 N41242 N41243 10
D41243 N41243 0 diode
R41244 N41243 N41244 10
D41244 N41244 0 diode
R41245 N41244 N41245 10
D41245 N41245 0 diode
R41246 N41245 N41246 10
D41246 N41246 0 diode
R41247 N41246 N41247 10
D41247 N41247 0 diode
R41248 N41247 N41248 10
D41248 N41248 0 diode
R41249 N41248 N41249 10
D41249 N41249 0 diode
R41250 N41249 N41250 10
D41250 N41250 0 diode
R41251 N41250 N41251 10
D41251 N41251 0 diode
R41252 N41251 N41252 10
D41252 N41252 0 diode
R41253 N41252 N41253 10
D41253 N41253 0 diode
R41254 N41253 N41254 10
D41254 N41254 0 diode
R41255 N41254 N41255 10
D41255 N41255 0 diode
R41256 N41255 N41256 10
D41256 N41256 0 diode
R41257 N41256 N41257 10
D41257 N41257 0 diode
R41258 N41257 N41258 10
D41258 N41258 0 diode
R41259 N41258 N41259 10
D41259 N41259 0 diode
R41260 N41259 N41260 10
D41260 N41260 0 diode
R41261 N41260 N41261 10
D41261 N41261 0 diode
R41262 N41261 N41262 10
D41262 N41262 0 diode
R41263 N41262 N41263 10
D41263 N41263 0 diode
R41264 N41263 N41264 10
D41264 N41264 0 diode
R41265 N41264 N41265 10
D41265 N41265 0 diode
R41266 N41265 N41266 10
D41266 N41266 0 diode
R41267 N41266 N41267 10
D41267 N41267 0 diode
R41268 N41267 N41268 10
D41268 N41268 0 diode
R41269 N41268 N41269 10
D41269 N41269 0 diode
R41270 N41269 N41270 10
D41270 N41270 0 diode
R41271 N41270 N41271 10
D41271 N41271 0 diode
R41272 N41271 N41272 10
D41272 N41272 0 diode
R41273 N41272 N41273 10
D41273 N41273 0 diode
R41274 N41273 N41274 10
D41274 N41274 0 diode
R41275 N41274 N41275 10
D41275 N41275 0 diode
R41276 N41275 N41276 10
D41276 N41276 0 diode
R41277 N41276 N41277 10
D41277 N41277 0 diode
R41278 N41277 N41278 10
D41278 N41278 0 diode
R41279 N41278 N41279 10
D41279 N41279 0 diode
R41280 N41279 N41280 10
D41280 N41280 0 diode
R41281 N41280 N41281 10
D41281 N41281 0 diode
R41282 N41281 N41282 10
D41282 N41282 0 diode
R41283 N41282 N41283 10
D41283 N41283 0 diode
R41284 N41283 N41284 10
D41284 N41284 0 diode
R41285 N41284 N41285 10
D41285 N41285 0 diode
R41286 N41285 N41286 10
D41286 N41286 0 diode
R41287 N41286 N41287 10
D41287 N41287 0 diode
R41288 N41287 N41288 10
D41288 N41288 0 diode
R41289 N41288 N41289 10
D41289 N41289 0 diode
R41290 N41289 N41290 10
D41290 N41290 0 diode
R41291 N41290 N41291 10
D41291 N41291 0 diode
R41292 N41291 N41292 10
D41292 N41292 0 diode
R41293 N41292 N41293 10
D41293 N41293 0 diode
R41294 N41293 N41294 10
D41294 N41294 0 diode
R41295 N41294 N41295 10
D41295 N41295 0 diode
R41296 N41295 N41296 10
D41296 N41296 0 diode
R41297 N41296 N41297 10
D41297 N41297 0 diode
R41298 N41297 N41298 10
D41298 N41298 0 diode
R41299 N41298 N41299 10
D41299 N41299 0 diode
R41300 N41299 N41300 10
D41300 N41300 0 diode
R41301 N41300 N41301 10
D41301 N41301 0 diode
R41302 N41301 N41302 10
D41302 N41302 0 diode
R41303 N41302 N41303 10
D41303 N41303 0 diode
R41304 N41303 N41304 10
D41304 N41304 0 diode
R41305 N41304 N41305 10
D41305 N41305 0 diode
R41306 N41305 N41306 10
D41306 N41306 0 diode
R41307 N41306 N41307 10
D41307 N41307 0 diode
R41308 N41307 N41308 10
D41308 N41308 0 diode
R41309 N41308 N41309 10
D41309 N41309 0 diode
R41310 N41309 N41310 10
D41310 N41310 0 diode
R41311 N41310 N41311 10
D41311 N41311 0 diode
R41312 N41311 N41312 10
D41312 N41312 0 diode
R41313 N41312 N41313 10
D41313 N41313 0 diode
R41314 N41313 N41314 10
D41314 N41314 0 diode
R41315 N41314 N41315 10
D41315 N41315 0 diode
R41316 N41315 N41316 10
D41316 N41316 0 diode
R41317 N41316 N41317 10
D41317 N41317 0 diode
R41318 N41317 N41318 10
D41318 N41318 0 diode
R41319 N41318 N41319 10
D41319 N41319 0 diode
R41320 N41319 N41320 10
D41320 N41320 0 diode
R41321 N41320 N41321 10
D41321 N41321 0 diode
R41322 N41321 N41322 10
D41322 N41322 0 diode
R41323 N41322 N41323 10
D41323 N41323 0 diode
R41324 N41323 N41324 10
D41324 N41324 0 diode
R41325 N41324 N41325 10
D41325 N41325 0 diode
R41326 N41325 N41326 10
D41326 N41326 0 diode
R41327 N41326 N41327 10
D41327 N41327 0 diode
R41328 N41327 N41328 10
D41328 N41328 0 diode
R41329 N41328 N41329 10
D41329 N41329 0 diode
R41330 N41329 N41330 10
D41330 N41330 0 diode
R41331 N41330 N41331 10
D41331 N41331 0 diode
R41332 N41331 N41332 10
D41332 N41332 0 diode
R41333 N41332 N41333 10
D41333 N41333 0 diode
R41334 N41333 N41334 10
D41334 N41334 0 diode
R41335 N41334 N41335 10
D41335 N41335 0 diode
R41336 N41335 N41336 10
D41336 N41336 0 diode
R41337 N41336 N41337 10
D41337 N41337 0 diode
R41338 N41337 N41338 10
D41338 N41338 0 diode
R41339 N41338 N41339 10
D41339 N41339 0 diode
R41340 N41339 N41340 10
D41340 N41340 0 diode
R41341 N41340 N41341 10
D41341 N41341 0 diode
R41342 N41341 N41342 10
D41342 N41342 0 diode
R41343 N41342 N41343 10
D41343 N41343 0 diode
R41344 N41343 N41344 10
D41344 N41344 0 diode
R41345 N41344 N41345 10
D41345 N41345 0 diode
R41346 N41345 N41346 10
D41346 N41346 0 diode
R41347 N41346 N41347 10
D41347 N41347 0 diode
R41348 N41347 N41348 10
D41348 N41348 0 diode
R41349 N41348 N41349 10
D41349 N41349 0 diode
R41350 N41349 N41350 10
D41350 N41350 0 diode
R41351 N41350 N41351 10
D41351 N41351 0 diode
R41352 N41351 N41352 10
D41352 N41352 0 diode
R41353 N41352 N41353 10
D41353 N41353 0 diode
R41354 N41353 N41354 10
D41354 N41354 0 diode
R41355 N41354 N41355 10
D41355 N41355 0 diode
R41356 N41355 N41356 10
D41356 N41356 0 diode
R41357 N41356 N41357 10
D41357 N41357 0 diode
R41358 N41357 N41358 10
D41358 N41358 0 diode
R41359 N41358 N41359 10
D41359 N41359 0 diode
R41360 N41359 N41360 10
D41360 N41360 0 diode
R41361 N41360 N41361 10
D41361 N41361 0 diode
R41362 N41361 N41362 10
D41362 N41362 0 diode
R41363 N41362 N41363 10
D41363 N41363 0 diode
R41364 N41363 N41364 10
D41364 N41364 0 diode
R41365 N41364 N41365 10
D41365 N41365 0 diode
R41366 N41365 N41366 10
D41366 N41366 0 diode
R41367 N41366 N41367 10
D41367 N41367 0 diode
R41368 N41367 N41368 10
D41368 N41368 0 diode
R41369 N41368 N41369 10
D41369 N41369 0 diode
R41370 N41369 N41370 10
D41370 N41370 0 diode
R41371 N41370 N41371 10
D41371 N41371 0 diode
R41372 N41371 N41372 10
D41372 N41372 0 diode
R41373 N41372 N41373 10
D41373 N41373 0 diode
R41374 N41373 N41374 10
D41374 N41374 0 diode
R41375 N41374 N41375 10
D41375 N41375 0 diode
R41376 N41375 N41376 10
D41376 N41376 0 diode
R41377 N41376 N41377 10
D41377 N41377 0 diode
R41378 N41377 N41378 10
D41378 N41378 0 diode
R41379 N41378 N41379 10
D41379 N41379 0 diode
R41380 N41379 N41380 10
D41380 N41380 0 diode
R41381 N41380 N41381 10
D41381 N41381 0 diode
R41382 N41381 N41382 10
D41382 N41382 0 diode
R41383 N41382 N41383 10
D41383 N41383 0 diode
R41384 N41383 N41384 10
D41384 N41384 0 diode
R41385 N41384 N41385 10
D41385 N41385 0 diode
R41386 N41385 N41386 10
D41386 N41386 0 diode
R41387 N41386 N41387 10
D41387 N41387 0 diode
R41388 N41387 N41388 10
D41388 N41388 0 diode
R41389 N41388 N41389 10
D41389 N41389 0 diode
R41390 N41389 N41390 10
D41390 N41390 0 diode
R41391 N41390 N41391 10
D41391 N41391 0 diode
R41392 N41391 N41392 10
D41392 N41392 0 diode
R41393 N41392 N41393 10
D41393 N41393 0 diode
R41394 N41393 N41394 10
D41394 N41394 0 diode
R41395 N41394 N41395 10
D41395 N41395 0 diode
R41396 N41395 N41396 10
D41396 N41396 0 diode
R41397 N41396 N41397 10
D41397 N41397 0 diode
R41398 N41397 N41398 10
D41398 N41398 0 diode
R41399 N41398 N41399 10
D41399 N41399 0 diode
R41400 N41399 N41400 10
D41400 N41400 0 diode
R41401 N41400 N41401 10
D41401 N41401 0 diode
R41402 N41401 N41402 10
D41402 N41402 0 diode
R41403 N41402 N41403 10
D41403 N41403 0 diode
R41404 N41403 N41404 10
D41404 N41404 0 diode
R41405 N41404 N41405 10
D41405 N41405 0 diode
R41406 N41405 N41406 10
D41406 N41406 0 diode
R41407 N41406 N41407 10
D41407 N41407 0 diode
R41408 N41407 N41408 10
D41408 N41408 0 diode
R41409 N41408 N41409 10
D41409 N41409 0 diode
R41410 N41409 N41410 10
D41410 N41410 0 diode
R41411 N41410 N41411 10
D41411 N41411 0 diode
R41412 N41411 N41412 10
D41412 N41412 0 diode
R41413 N41412 N41413 10
D41413 N41413 0 diode
R41414 N41413 N41414 10
D41414 N41414 0 diode
R41415 N41414 N41415 10
D41415 N41415 0 diode
R41416 N41415 N41416 10
D41416 N41416 0 diode
R41417 N41416 N41417 10
D41417 N41417 0 diode
R41418 N41417 N41418 10
D41418 N41418 0 diode
R41419 N41418 N41419 10
D41419 N41419 0 diode
R41420 N41419 N41420 10
D41420 N41420 0 diode
R41421 N41420 N41421 10
D41421 N41421 0 diode
R41422 N41421 N41422 10
D41422 N41422 0 diode
R41423 N41422 N41423 10
D41423 N41423 0 diode
R41424 N41423 N41424 10
D41424 N41424 0 diode
R41425 N41424 N41425 10
D41425 N41425 0 diode
R41426 N41425 N41426 10
D41426 N41426 0 diode
R41427 N41426 N41427 10
D41427 N41427 0 diode
R41428 N41427 N41428 10
D41428 N41428 0 diode
R41429 N41428 N41429 10
D41429 N41429 0 diode
R41430 N41429 N41430 10
D41430 N41430 0 diode
R41431 N41430 N41431 10
D41431 N41431 0 diode
R41432 N41431 N41432 10
D41432 N41432 0 diode
R41433 N41432 N41433 10
D41433 N41433 0 diode
R41434 N41433 N41434 10
D41434 N41434 0 diode
R41435 N41434 N41435 10
D41435 N41435 0 diode
R41436 N41435 N41436 10
D41436 N41436 0 diode
R41437 N41436 N41437 10
D41437 N41437 0 diode
R41438 N41437 N41438 10
D41438 N41438 0 diode
R41439 N41438 N41439 10
D41439 N41439 0 diode
R41440 N41439 N41440 10
D41440 N41440 0 diode
R41441 N41440 N41441 10
D41441 N41441 0 diode
R41442 N41441 N41442 10
D41442 N41442 0 diode
R41443 N41442 N41443 10
D41443 N41443 0 diode
R41444 N41443 N41444 10
D41444 N41444 0 diode
R41445 N41444 N41445 10
D41445 N41445 0 diode
R41446 N41445 N41446 10
D41446 N41446 0 diode
R41447 N41446 N41447 10
D41447 N41447 0 diode
R41448 N41447 N41448 10
D41448 N41448 0 diode
R41449 N41448 N41449 10
D41449 N41449 0 diode
R41450 N41449 N41450 10
D41450 N41450 0 diode
R41451 N41450 N41451 10
D41451 N41451 0 diode
R41452 N41451 N41452 10
D41452 N41452 0 diode
R41453 N41452 N41453 10
D41453 N41453 0 diode
R41454 N41453 N41454 10
D41454 N41454 0 diode
R41455 N41454 N41455 10
D41455 N41455 0 diode
R41456 N41455 N41456 10
D41456 N41456 0 diode
R41457 N41456 N41457 10
D41457 N41457 0 diode
R41458 N41457 N41458 10
D41458 N41458 0 diode
R41459 N41458 N41459 10
D41459 N41459 0 diode
R41460 N41459 N41460 10
D41460 N41460 0 diode
R41461 N41460 N41461 10
D41461 N41461 0 diode
R41462 N41461 N41462 10
D41462 N41462 0 diode
R41463 N41462 N41463 10
D41463 N41463 0 diode
R41464 N41463 N41464 10
D41464 N41464 0 diode
R41465 N41464 N41465 10
D41465 N41465 0 diode
R41466 N41465 N41466 10
D41466 N41466 0 diode
R41467 N41466 N41467 10
D41467 N41467 0 diode
R41468 N41467 N41468 10
D41468 N41468 0 diode
R41469 N41468 N41469 10
D41469 N41469 0 diode
R41470 N41469 N41470 10
D41470 N41470 0 diode
R41471 N41470 N41471 10
D41471 N41471 0 diode
R41472 N41471 N41472 10
D41472 N41472 0 diode
R41473 N41472 N41473 10
D41473 N41473 0 diode
R41474 N41473 N41474 10
D41474 N41474 0 diode
R41475 N41474 N41475 10
D41475 N41475 0 diode
R41476 N41475 N41476 10
D41476 N41476 0 diode
R41477 N41476 N41477 10
D41477 N41477 0 diode
R41478 N41477 N41478 10
D41478 N41478 0 diode
R41479 N41478 N41479 10
D41479 N41479 0 diode
R41480 N41479 N41480 10
D41480 N41480 0 diode
R41481 N41480 N41481 10
D41481 N41481 0 diode
R41482 N41481 N41482 10
D41482 N41482 0 diode
R41483 N41482 N41483 10
D41483 N41483 0 diode
R41484 N41483 N41484 10
D41484 N41484 0 diode
R41485 N41484 N41485 10
D41485 N41485 0 diode
R41486 N41485 N41486 10
D41486 N41486 0 diode
R41487 N41486 N41487 10
D41487 N41487 0 diode
R41488 N41487 N41488 10
D41488 N41488 0 diode
R41489 N41488 N41489 10
D41489 N41489 0 diode
R41490 N41489 N41490 10
D41490 N41490 0 diode
R41491 N41490 N41491 10
D41491 N41491 0 diode
R41492 N41491 N41492 10
D41492 N41492 0 diode
R41493 N41492 N41493 10
D41493 N41493 0 diode
R41494 N41493 N41494 10
D41494 N41494 0 diode
R41495 N41494 N41495 10
D41495 N41495 0 diode
R41496 N41495 N41496 10
D41496 N41496 0 diode
R41497 N41496 N41497 10
D41497 N41497 0 diode
R41498 N41497 N41498 10
D41498 N41498 0 diode
R41499 N41498 N41499 10
D41499 N41499 0 diode
R41500 N41499 N41500 10
D41500 N41500 0 diode
R41501 N41500 N41501 10
D41501 N41501 0 diode
R41502 N41501 N41502 10
D41502 N41502 0 diode
R41503 N41502 N41503 10
D41503 N41503 0 diode
R41504 N41503 N41504 10
D41504 N41504 0 diode
R41505 N41504 N41505 10
D41505 N41505 0 diode
R41506 N41505 N41506 10
D41506 N41506 0 diode
R41507 N41506 N41507 10
D41507 N41507 0 diode
R41508 N41507 N41508 10
D41508 N41508 0 diode
R41509 N41508 N41509 10
D41509 N41509 0 diode
R41510 N41509 N41510 10
D41510 N41510 0 diode
R41511 N41510 N41511 10
D41511 N41511 0 diode
R41512 N41511 N41512 10
D41512 N41512 0 diode
R41513 N41512 N41513 10
D41513 N41513 0 diode
R41514 N41513 N41514 10
D41514 N41514 0 diode
R41515 N41514 N41515 10
D41515 N41515 0 diode
R41516 N41515 N41516 10
D41516 N41516 0 diode
R41517 N41516 N41517 10
D41517 N41517 0 diode
R41518 N41517 N41518 10
D41518 N41518 0 diode
R41519 N41518 N41519 10
D41519 N41519 0 diode
R41520 N41519 N41520 10
D41520 N41520 0 diode
R41521 N41520 N41521 10
D41521 N41521 0 diode
R41522 N41521 N41522 10
D41522 N41522 0 diode
R41523 N41522 N41523 10
D41523 N41523 0 diode
R41524 N41523 N41524 10
D41524 N41524 0 diode
R41525 N41524 N41525 10
D41525 N41525 0 diode
R41526 N41525 N41526 10
D41526 N41526 0 diode
R41527 N41526 N41527 10
D41527 N41527 0 diode
R41528 N41527 N41528 10
D41528 N41528 0 diode
R41529 N41528 N41529 10
D41529 N41529 0 diode
R41530 N41529 N41530 10
D41530 N41530 0 diode
R41531 N41530 N41531 10
D41531 N41531 0 diode
R41532 N41531 N41532 10
D41532 N41532 0 diode
R41533 N41532 N41533 10
D41533 N41533 0 diode
R41534 N41533 N41534 10
D41534 N41534 0 diode
R41535 N41534 N41535 10
D41535 N41535 0 diode
R41536 N41535 N41536 10
D41536 N41536 0 diode
R41537 N41536 N41537 10
D41537 N41537 0 diode
R41538 N41537 N41538 10
D41538 N41538 0 diode
R41539 N41538 N41539 10
D41539 N41539 0 diode
R41540 N41539 N41540 10
D41540 N41540 0 diode
R41541 N41540 N41541 10
D41541 N41541 0 diode
R41542 N41541 N41542 10
D41542 N41542 0 diode
R41543 N41542 N41543 10
D41543 N41543 0 diode
R41544 N41543 N41544 10
D41544 N41544 0 diode
R41545 N41544 N41545 10
D41545 N41545 0 diode
R41546 N41545 N41546 10
D41546 N41546 0 diode
R41547 N41546 N41547 10
D41547 N41547 0 diode
R41548 N41547 N41548 10
D41548 N41548 0 diode
R41549 N41548 N41549 10
D41549 N41549 0 diode
R41550 N41549 N41550 10
D41550 N41550 0 diode
R41551 N41550 N41551 10
D41551 N41551 0 diode
R41552 N41551 N41552 10
D41552 N41552 0 diode
R41553 N41552 N41553 10
D41553 N41553 0 diode
R41554 N41553 N41554 10
D41554 N41554 0 diode
R41555 N41554 N41555 10
D41555 N41555 0 diode
R41556 N41555 N41556 10
D41556 N41556 0 diode
R41557 N41556 N41557 10
D41557 N41557 0 diode
R41558 N41557 N41558 10
D41558 N41558 0 diode
R41559 N41558 N41559 10
D41559 N41559 0 diode
R41560 N41559 N41560 10
D41560 N41560 0 diode
R41561 N41560 N41561 10
D41561 N41561 0 diode
R41562 N41561 N41562 10
D41562 N41562 0 diode
R41563 N41562 N41563 10
D41563 N41563 0 diode
R41564 N41563 N41564 10
D41564 N41564 0 diode
R41565 N41564 N41565 10
D41565 N41565 0 diode
R41566 N41565 N41566 10
D41566 N41566 0 diode
R41567 N41566 N41567 10
D41567 N41567 0 diode
R41568 N41567 N41568 10
D41568 N41568 0 diode
R41569 N41568 N41569 10
D41569 N41569 0 diode
R41570 N41569 N41570 10
D41570 N41570 0 diode
R41571 N41570 N41571 10
D41571 N41571 0 diode
R41572 N41571 N41572 10
D41572 N41572 0 diode
R41573 N41572 N41573 10
D41573 N41573 0 diode
R41574 N41573 N41574 10
D41574 N41574 0 diode
R41575 N41574 N41575 10
D41575 N41575 0 diode
R41576 N41575 N41576 10
D41576 N41576 0 diode
R41577 N41576 N41577 10
D41577 N41577 0 diode
R41578 N41577 N41578 10
D41578 N41578 0 diode
R41579 N41578 N41579 10
D41579 N41579 0 diode
R41580 N41579 N41580 10
D41580 N41580 0 diode
R41581 N41580 N41581 10
D41581 N41581 0 diode
R41582 N41581 N41582 10
D41582 N41582 0 diode
R41583 N41582 N41583 10
D41583 N41583 0 diode
R41584 N41583 N41584 10
D41584 N41584 0 diode
R41585 N41584 N41585 10
D41585 N41585 0 diode
R41586 N41585 N41586 10
D41586 N41586 0 diode
R41587 N41586 N41587 10
D41587 N41587 0 diode
R41588 N41587 N41588 10
D41588 N41588 0 diode
R41589 N41588 N41589 10
D41589 N41589 0 diode
R41590 N41589 N41590 10
D41590 N41590 0 diode
R41591 N41590 N41591 10
D41591 N41591 0 diode
R41592 N41591 N41592 10
D41592 N41592 0 diode
R41593 N41592 N41593 10
D41593 N41593 0 diode
R41594 N41593 N41594 10
D41594 N41594 0 diode
R41595 N41594 N41595 10
D41595 N41595 0 diode
R41596 N41595 N41596 10
D41596 N41596 0 diode
R41597 N41596 N41597 10
D41597 N41597 0 diode
R41598 N41597 N41598 10
D41598 N41598 0 diode
R41599 N41598 N41599 10
D41599 N41599 0 diode
R41600 N41599 N41600 10
D41600 N41600 0 diode
R41601 N41600 N41601 10
D41601 N41601 0 diode
R41602 N41601 N41602 10
D41602 N41602 0 diode
R41603 N41602 N41603 10
D41603 N41603 0 diode
R41604 N41603 N41604 10
D41604 N41604 0 diode
R41605 N41604 N41605 10
D41605 N41605 0 diode
R41606 N41605 N41606 10
D41606 N41606 0 diode
R41607 N41606 N41607 10
D41607 N41607 0 diode
R41608 N41607 N41608 10
D41608 N41608 0 diode
R41609 N41608 N41609 10
D41609 N41609 0 diode
R41610 N41609 N41610 10
D41610 N41610 0 diode
R41611 N41610 N41611 10
D41611 N41611 0 diode
R41612 N41611 N41612 10
D41612 N41612 0 diode
R41613 N41612 N41613 10
D41613 N41613 0 diode
R41614 N41613 N41614 10
D41614 N41614 0 diode
R41615 N41614 N41615 10
D41615 N41615 0 diode
R41616 N41615 N41616 10
D41616 N41616 0 diode
R41617 N41616 N41617 10
D41617 N41617 0 diode
R41618 N41617 N41618 10
D41618 N41618 0 diode
R41619 N41618 N41619 10
D41619 N41619 0 diode
R41620 N41619 N41620 10
D41620 N41620 0 diode
R41621 N41620 N41621 10
D41621 N41621 0 diode
R41622 N41621 N41622 10
D41622 N41622 0 diode
R41623 N41622 N41623 10
D41623 N41623 0 diode
R41624 N41623 N41624 10
D41624 N41624 0 diode
R41625 N41624 N41625 10
D41625 N41625 0 diode
R41626 N41625 N41626 10
D41626 N41626 0 diode
R41627 N41626 N41627 10
D41627 N41627 0 diode
R41628 N41627 N41628 10
D41628 N41628 0 diode
R41629 N41628 N41629 10
D41629 N41629 0 diode
R41630 N41629 N41630 10
D41630 N41630 0 diode
R41631 N41630 N41631 10
D41631 N41631 0 diode
R41632 N41631 N41632 10
D41632 N41632 0 diode
R41633 N41632 N41633 10
D41633 N41633 0 diode
R41634 N41633 N41634 10
D41634 N41634 0 diode
R41635 N41634 N41635 10
D41635 N41635 0 diode
R41636 N41635 N41636 10
D41636 N41636 0 diode
R41637 N41636 N41637 10
D41637 N41637 0 diode
R41638 N41637 N41638 10
D41638 N41638 0 diode
R41639 N41638 N41639 10
D41639 N41639 0 diode
R41640 N41639 N41640 10
D41640 N41640 0 diode
R41641 N41640 N41641 10
D41641 N41641 0 diode
R41642 N41641 N41642 10
D41642 N41642 0 diode
R41643 N41642 N41643 10
D41643 N41643 0 diode
R41644 N41643 N41644 10
D41644 N41644 0 diode
R41645 N41644 N41645 10
D41645 N41645 0 diode
R41646 N41645 N41646 10
D41646 N41646 0 diode
R41647 N41646 N41647 10
D41647 N41647 0 diode
R41648 N41647 N41648 10
D41648 N41648 0 diode
R41649 N41648 N41649 10
D41649 N41649 0 diode
R41650 N41649 N41650 10
D41650 N41650 0 diode
R41651 N41650 N41651 10
D41651 N41651 0 diode
R41652 N41651 N41652 10
D41652 N41652 0 diode
R41653 N41652 N41653 10
D41653 N41653 0 diode
R41654 N41653 N41654 10
D41654 N41654 0 diode
R41655 N41654 N41655 10
D41655 N41655 0 diode
R41656 N41655 N41656 10
D41656 N41656 0 diode
R41657 N41656 N41657 10
D41657 N41657 0 diode
R41658 N41657 N41658 10
D41658 N41658 0 diode
R41659 N41658 N41659 10
D41659 N41659 0 diode
R41660 N41659 N41660 10
D41660 N41660 0 diode
R41661 N41660 N41661 10
D41661 N41661 0 diode
R41662 N41661 N41662 10
D41662 N41662 0 diode
R41663 N41662 N41663 10
D41663 N41663 0 diode
R41664 N41663 N41664 10
D41664 N41664 0 diode
R41665 N41664 N41665 10
D41665 N41665 0 diode
R41666 N41665 N41666 10
D41666 N41666 0 diode
R41667 N41666 N41667 10
D41667 N41667 0 diode
R41668 N41667 N41668 10
D41668 N41668 0 diode
R41669 N41668 N41669 10
D41669 N41669 0 diode
R41670 N41669 N41670 10
D41670 N41670 0 diode
R41671 N41670 N41671 10
D41671 N41671 0 diode
R41672 N41671 N41672 10
D41672 N41672 0 diode
R41673 N41672 N41673 10
D41673 N41673 0 diode
R41674 N41673 N41674 10
D41674 N41674 0 diode
R41675 N41674 N41675 10
D41675 N41675 0 diode
R41676 N41675 N41676 10
D41676 N41676 0 diode
R41677 N41676 N41677 10
D41677 N41677 0 diode
R41678 N41677 N41678 10
D41678 N41678 0 diode
R41679 N41678 N41679 10
D41679 N41679 0 diode
R41680 N41679 N41680 10
D41680 N41680 0 diode
R41681 N41680 N41681 10
D41681 N41681 0 diode
R41682 N41681 N41682 10
D41682 N41682 0 diode
R41683 N41682 N41683 10
D41683 N41683 0 diode
R41684 N41683 N41684 10
D41684 N41684 0 diode
R41685 N41684 N41685 10
D41685 N41685 0 diode
R41686 N41685 N41686 10
D41686 N41686 0 diode
R41687 N41686 N41687 10
D41687 N41687 0 diode
R41688 N41687 N41688 10
D41688 N41688 0 diode
R41689 N41688 N41689 10
D41689 N41689 0 diode
R41690 N41689 N41690 10
D41690 N41690 0 diode
R41691 N41690 N41691 10
D41691 N41691 0 diode
R41692 N41691 N41692 10
D41692 N41692 0 diode
R41693 N41692 N41693 10
D41693 N41693 0 diode
R41694 N41693 N41694 10
D41694 N41694 0 diode
R41695 N41694 N41695 10
D41695 N41695 0 diode
R41696 N41695 N41696 10
D41696 N41696 0 diode
R41697 N41696 N41697 10
D41697 N41697 0 diode
R41698 N41697 N41698 10
D41698 N41698 0 diode
R41699 N41698 N41699 10
D41699 N41699 0 diode
R41700 N41699 N41700 10
D41700 N41700 0 diode
R41701 N41700 N41701 10
D41701 N41701 0 diode
R41702 N41701 N41702 10
D41702 N41702 0 diode
R41703 N41702 N41703 10
D41703 N41703 0 diode
R41704 N41703 N41704 10
D41704 N41704 0 diode
R41705 N41704 N41705 10
D41705 N41705 0 diode
R41706 N41705 N41706 10
D41706 N41706 0 diode
R41707 N41706 N41707 10
D41707 N41707 0 diode
R41708 N41707 N41708 10
D41708 N41708 0 diode
R41709 N41708 N41709 10
D41709 N41709 0 diode
R41710 N41709 N41710 10
D41710 N41710 0 diode
R41711 N41710 N41711 10
D41711 N41711 0 diode
R41712 N41711 N41712 10
D41712 N41712 0 diode
R41713 N41712 N41713 10
D41713 N41713 0 diode
R41714 N41713 N41714 10
D41714 N41714 0 diode
R41715 N41714 N41715 10
D41715 N41715 0 diode
R41716 N41715 N41716 10
D41716 N41716 0 diode
R41717 N41716 N41717 10
D41717 N41717 0 diode
R41718 N41717 N41718 10
D41718 N41718 0 diode
R41719 N41718 N41719 10
D41719 N41719 0 diode
R41720 N41719 N41720 10
D41720 N41720 0 diode
R41721 N41720 N41721 10
D41721 N41721 0 diode
R41722 N41721 N41722 10
D41722 N41722 0 diode
R41723 N41722 N41723 10
D41723 N41723 0 diode
R41724 N41723 N41724 10
D41724 N41724 0 diode
R41725 N41724 N41725 10
D41725 N41725 0 diode
R41726 N41725 N41726 10
D41726 N41726 0 diode
R41727 N41726 N41727 10
D41727 N41727 0 diode
R41728 N41727 N41728 10
D41728 N41728 0 diode
R41729 N41728 N41729 10
D41729 N41729 0 diode
R41730 N41729 N41730 10
D41730 N41730 0 diode
R41731 N41730 N41731 10
D41731 N41731 0 diode
R41732 N41731 N41732 10
D41732 N41732 0 diode
R41733 N41732 N41733 10
D41733 N41733 0 diode
R41734 N41733 N41734 10
D41734 N41734 0 diode
R41735 N41734 N41735 10
D41735 N41735 0 diode
R41736 N41735 N41736 10
D41736 N41736 0 diode
R41737 N41736 N41737 10
D41737 N41737 0 diode
R41738 N41737 N41738 10
D41738 N41738 0 diode
R41739 N41738 N41739 10
D41739 N41739 0 diode
R41740 N41739 N41740 10
D41740 N41740 0 diode
R41741 N41740 N41741 10
D41741 N41741 0 diode
R41742 N41741 N41742 10
D41742 N41742 0 diode
R41743 N41742 N41743 10
D41743 N41743 0 diode
R41744 N41743 N41744 10
D41744 N41744 0 diode
R41745 N41744 N41745 10
D41745 N41745 0 diode
R41746 N41745 N41746 10
D41746 N41746 0 diode
R41747 N41746 N41747 10
D41747 N41747 0 diode
R41748 N41747 N41748 10
D41748 N41748 0 diode
R41749 N41748 N41749 10
D41749 N41749 0 diode
R41750 N41749 N41750 10
D41750 N41750 0 diode
R41751 N41750 N41751 10
D41751 N41751 0 diode
R41752 N41751 N41752 10
D41752 N41752 0 diode
R41753 N41752 N41753 10
D41753 N41753 0 diode
R41754 N41753 N41754 10
D41754 N41754 0 diode
R41755 N41754 N41755 10
D41755 N41755 0 diode
R41756 N41755 N41756 10
D41756 N41756 0 diode
R41757 N41756 N41757 10
D41757 N41757 0 diode
R41758 N41757 N41758 10
D41758 N41758 0 diode
R41759 N41758 N41759 10
D41759 N41759 0 diode
R41760 N41759 N41760 10
D41760 N41760 0 diode
R41761 N41760 N41761 10
D41761 N41761 0 diode
R41762 N41761 N41762 10
D41762 N41762 0 diode
R41763 N41762 N41763 10
D41763 N41763 0 diode
R41764 N41763 N41764 10
D41764 N41764 0 diode
R41765 N41764 N41765 10
D41765 N41765 0 diode
R41766 N41765 N41766 10
D41766 N41766 0 diode
R41767 N41766 N41767 10
D41767 N41767 0 diode
R41768 N41767 N41768 10
D41768 N41768 0 diode
R41769 N41768 N41769 10
D41769 N41769 0 diode
R41770 N41769 N41770 10
D41770 N41770 0 diode
R41771 N41770 N41771 10
D41771 N41771 0 diode
R41772 N41771 N41772 10
D41772 N41772 0 diode
R41773 N41772 N41773 10
D41773 N41773 0 diode
R41774 N41773 N41774 10
D41774 N41774 0 diode
R41775 N41774 N41775 10
D41775 N41775 0 diode
R41776 N41775 N41776 10
D41776 N41776 0 diode
R41777 N41776 N41777 10
D41777 N41777 0 diode
R41778 N41777 N41778 10
D41778 N41778 0 diode
R41779 N41778 N41779 10
D41779 N41779 0 diode
R41780 N41779 N41780 10
D41780 N41780 0 diode
R41781 N41780 N41781 10
D41781 N41781 0 diode
R41782 N41781 N41782 10
D41782 N41782 0 diode
R41783 N41782 N41783 10
D41783 N41783 0 diode
R41784 N41783 N41784 10
D41784 N41784 0 diode
R41785 N41784 N41785 10
D41785 N41785 0 diode
R41786 N41785 N41786 10
D41786 N41786 0 diode
R41787 N41786 N41787 10
D41787 N41787 0 diode
R41788 N41787 N41788 10
D41788 N41788 0 diode
R41789 N41788 N41789 10
D41789 N41789 0 diode
R41790 N41789 N41790 10
D41790 N41790 0 diode
R41791 N41790 N41791 10
D41791 N41791 0 diode
R41792 N41791 N41792 10
D41792 N41792 0 diode
R41793 N41792 N41793 10
D41793 N41793 0 diode
R41794 N41793 N41794 10
D41794 N41794 0 diode
R41795 N41794 N41795 10
D41795 N41795 0 diode
R41796 N41795 N41796 10
D41796 N41796 0 diode
R41797 N41796 N41797 10
D41797 N41797 0 diode
R41798 N41797 N41798 10
D41798 N41798 0 diode
R41799 N41798 N41799 10
D41799 N41799 0 diode
R41800 N41799 N41800 10
D41800 N41800 0 diode
R41801 N41800 N41801 10
D41801 N41801 0 diode
R41802 N41801 N41802 10
D41802 N41802 0 diode
R41803 N41802 N41803 10
D41803 N41803 0 diode
R41804 N41803 N41804 10
D41804 N41804 0 diode
R41805 N41804 N41805 10
D41805 N41805 0 diode
R41806 N41805 N41806 10
D41806 N41806 0 diode
R41807 N41806 N41807 10
D41807 N41807 0 diode
R41808 N41807 N41808 10
D41808 N41808 0 diode
R41809 N41808 N41809 10
D41809 N41809 0 diode
R41810 N41809 N41810 10
D41810 N41810 0 diode
R41811 N41810 N41811 10
D41811 N41811 0 diode
R41812 N41811 N41812 10
D41812 N41812 0 diode
R41813 N41812 N41813 10
D41813 N41813 0 diode
R41814 N41813 N41814 10
D41814 N41814 0 diode
R41815 N41814 N41815 10
D41815 N41815 0 diode
R41816 N41815 N41816 10
D41816 N41816 0 diode
R41817 N41816 N41817 10
D41817 N41817 0 diode
R41818 N41817 N41818 10
D41818 N41818 0 diode
R41819 N41818 N41819 10
D41819 N41819 0 diode
R41820 N41819 N41820 10
D41820 N41820 0 diode
R41821 N41820 N41821 10
D41821 N41821 0 diode
R41822 N41821 N41822 10
D41822 N41822 0 diode
R41823 N41822 N41823 10
D41823 N41823 0 diode
R41824 N41823 N41824 10
D41824 N41824 0 diode
R41825 N41824 N41825 10
D41825 N41825 0 diode
R41826 N41825 N41826 10
D41826 N41826 0 diode
R41827 N41826 N41827 10
D41827 N41827 0 diode
R41828 N41827 N41828 10
D41828 N41828 0 diode
R41829 N41828 N41829 10
D41829 N41829 0 diode
R41830 N41829 N41830 10
D41830 N41830 0 diode
R41831 N41830 N41831 10
D41831 N41831 0 diode
R41832 N41831 N41832 10
D41832 N41832 0 diode
R41833 N41832 N41833 10
D41833 N41833 0 diode
R41834 N41833 N41834 10
D41834 N41834 0 diode
R41835 N41834 N41835 10
D41835 N41835 0 diode
R41836 N41835 N41836 10
D41836 N41836 0 diode
R41837 N41836 N41837 10
D41837 N41837 0 diode
R41838 N41837 N41838 10
D41838 N41838 0 diode
R41839 N41838 N41839 10
D41839 N41839 0 diode
R41840 N41839 N41840 10
D41840 N41840 0 diode
R41841 N41840 N41841 10
D41841 N41841 0 diode
R41842 N41841 N41842 10
D41842 N41842 0 diode
R41843 N41842 N41843 10
D41843 N41843 0 diode
R41844 N41843 N41844 10
D41844 N41844 0 diode
R41845 N41844 N41845 10
D41845 N41845 0 diode
R41846 N41845 N41846 10
D41846 N41846 0 diode
R41847 N41846 N41847 10
D41847 N41847 0 diode
R41848 N41847 N41848 10
D41848 N41848 0 diode
R41849 N41848 N41849 10
D41849 N41849 0 diode
R41850 N41849 N41850 10
D41850 N41850 0 diode
R41851 N41850 N41851 10
D41851 N41851 0 diode
R41852 N41851 N41852 10
D41852 N41852 0 diode
R41853 N41852 N41853 10
D41853 N41853 0 diode
R41854 N41853 N41854 10
D41854 N41854 0 diode
R41855 N41854 N41855 10
D41855 N41855 0 diode
R41856 N41855 N41856 10
D41856 N41856 0 diode
R41857 N41856 N41857 10
D41857 N41857 0 diode
R41858 N41857 N41858 10
D41858 N41858 0 diode
R41859 N41858 N41859 10
D41859 N41859 0 diode
R41860 N41859 N41860 10
D41860 N41860 0 diode
R41861 N41860 N41861 10
D41861 N41861 0 diode
R41862 N41861 N41862 10
D41862 N41862 0 diode
R41863 N41862 N41863 10
D41863 N41863 0 diode
R41864 N41863 N41864 10
D41864 N41864 0 diode
R41865 N41864 N41865 10
D41865 N41865 0 diode
R41866 N41865 N41866 10
D41866 N41866 0 diode
R41867 N41866 N41867 10
D41867 N41867 0 diode
R41868 N41867 N41868 10
D41868 N41868 0 diode
R41869 N41868 N41869 10
D41869 N41869 0 diode
R41870 N41869 N41870 10
D41870 N41870 0 diode
R41871 N41870 N41871 10
D41871 N41871 0 diode
R41872 N41871 N41872 10
D41872 N41872 0 diode
R41873 N41872 N41873 10
D41873 N41873 0 diode
R41874 N41873 N41874 10
D41874 N41874 0 diode
R41875 N41874 N41875 10
D41875 N41875 0 diode
R41876 N41875 N41876 10
D41876 N41876 0 diode
R41877 N41876 N41877 10
D41877 N41877 0 diode
R41878 N41877 N41878 10
D41878 N41878 0 diode
R41879 N41878 N41879 10
D41879 N41879 0 diode
R41880 N41879 N41880 10
D41880 N41880 0 diode
R41881 N41880 N41881 10
D41881 N41881 0 diode
R41882 N41881 N41882 10
D41882 N41882 0 diode
R41883 N41882 N41883 10
D41883 N41883 0 diode
R41884 N41883 N41884 10
D41884 N41884 0 diode
R41885 N41884 N41885 10
D41885 N41885 0 diode
R41886 N41885 N41886 10
D41886 N41886 0 diode
R41887 N41886 N41887 10
D41887 N41887 0 diode
R41888 N41887 N41888 10
D41888 N41888 0 diode
R41889 N41888 N41889 10
D41889 N41889 0 diode
R41890 N41889 N41890 10
D41890 N41890 0 diode
R41891 N41890 N41891 10
D41891 N41891 0 diode
R41892 N41891 N41892 10
D41892 N41892 0 diode
R41893 N41892 N41893 10
D41893 N41893 0 diode
R41894 N41893 N41894 10
D41894 N41894 0 diode
R41895 N41894 N41895 10
D41895 N41895 0 diode
R41896 N41895 N41896 10
D41896 N41896 0 diode
R41897 N41896 N41897 10
D41897 N41897 0 diode
R41898 N41897 N41898 10
D41898 N41898 0 diode
R41899 N41898 N41899 10
D41899 N41899 0 diode
R41900 N41899 N41900 10
D41900 N41900 0 diode
R41901 N41900 N41901 10
D41901 N41901 0 diode
R41902 N41901 N41902 10
D41902 N41902 0 diode
R41903 N41902 N41903 10
D41903 N41903 0 diode
R41904 N41903 N41904 10
D41904 N41904 0 diode
R41905 N41904 N41905 10
D41905 N41905 0 diode
R41906 N41905 N41906 10
D41906 N41906 0 diode
R41907 N41906 N41907 10
D41907 N41907 0 diode
R41908 N41907 N41908 10
D41908 N41908 0 diode
R41909 N41908 N41909 10
D41909 N41909 0 diode
R41910 N41909 N41910 10
D41910 N41910 0 diode
R41911 N41910 N41911 10
D41911 N41911 0 diode
R41912 N41911 N41912 10
D41912 N41912 0 diode
R41913 N41912 N41913 10
D41913 N41913 0 diode
R41914 N41913 N41914 10
D41914 N41914 0 diode
R41915 N41914 N41915 10
D41915 N41915 0 diode
R41916 N41915 N41916 10
D41916 N41916 0 diode
R41917 N41916 N41917 10
D41917 N41917 0 diode
R41918 N41917 N41918 10
D41918 N41918 0 diode
R41919 N41918 N41919 10
D41919 N41919 0 diode
R41920 N41919 N41920 10
D41920 N41920 0 diode
R41921 N41920 N41921 10
D41921 N41921 0 diode
R41922 N41921 N41922 10
D41922 N41922 0 diode
R41923 N41922 N41923 10
D41923 N41923 0 diode
R41924 N41923 N41924 10
D41924 N41924 0 diode
R41925 N41924 N41925 10
D41925 N41925 0 diode
R41926 N41925 N41926 10
D41926 N41926 0 diode
R41927 N41926 N41927 10
D41927 N41927 0 diode
R41928 N41927 N41928 10
D41928 N41928 0 diode
R41929 N41928 N41929 10
D41929 N41929 0 diode
R41930 N41929 N41930 10
D41930 N41930 0 diode
R41931 N41930 N41931 10
D41931 N41931 0 diode
R41932 N41931 N41932 10
D41932 N41932 0 diode
R41933 N41932 N41933 10
D41933 N41933 0 diode
R41934 N41933 N41934 10
D41934 N41934 0 diode
R41935 N41934 N41935 10
D41935 N41935 0 diode
R41936 N41935 N41936 10
D41936 N41936 0 diode
R41937 N41936 N41937 10
D41937 N41937 0 diode
R41938 N41937 N41938 10
D41938 N41938 0 diode
R41939 N41938 N41939 10
D41939 N41939 0 diode
R41940 N41939 N41940 10
D41940 N41940 0 diode
R41941 N41940 N41941 10
D41941 N41941 0 diode
R41942 N41941 N41942 10
D41942 N41942 0 diode
R41943 N41942 N41943 10
D41943 N41943 0 diode
R41944 N41943 N41944 10
D41944 N41944 0 diode
R41945 N41944 N41945 10
D41945 N41945 0 diode
R41946 N41945 N41946 10
D41946 N41946 0 diode
R41947 N41946 N41947 10
D41947 N41947 0 diode
R41948 N41947 N41948 10
D41948 N41948 0 diode
R41949 N41948 N41949 10
D41949 N41949 0 diode
R41950 N41949 N41950 10
D41950 N41950 0 diode
R41951 N41950 N41951 10
D41951 N41951 0 diode
R41952 N41951 N41952 10
D41952 N41952 0 diode
R41953 N41952 N41953 10
D41953 N41953 0 diode
R41954 N41953 N41954 10
D41954 N41954 0 diode
R41955 N41954 N41955 10
D41955 N41955 0 diode
R41956 N41955 N41956 10
D41956 N41956 0 diode
R41957 N41956 N41957 10
D41957 N41957 0 diode
R41958 N41957 N41958 10
D41958 N41958 0 diode
R41959 N41958 N41959 10
D41959 N41959 0 diode
R41960 N41959 N41960 10
D41960 N41960 0 diode
R41961 N41960 N41961 10
D41961 N41961 0 diode
R41962 N41961 N41962 10
D41962 N41962 0 diode
R41963 N41962 N41963 10
D41963 N41963 0 diode
R41964 N41963 N41964 10
D41964 N41964 0 diode
R41965 N41964 N41965 10
D41965 N41965 0 diode
R41966 N41965 N41966 10
D41966 N41966 0 diode
R41967 N41966 N41967 10
D41967 N41967 0 diode
R41968 N41967 N41968 10
D41968 N41968 0 diode
R41969 N41968 N41969 10
D41969 N41969 0 diode
R41970 N41969 N41970 10
D41970 N41970 0 diode
R41971 N41970 N41971 10
D41971 N41971 0 diode
R41972 N41971 N41972 10
D41972 N41972 0 diode
R41973 N41972 N41973 10
D41973 N41973 0 diode
R41974 N41973 N41974 10
D41974 N41974 0 diode
R41975 N41974 N41975 10
D41975 N41975 0 diode
R41976 N41975 N41976 10
D41976 N41976 0 diode
R41977 N41976 N41977 10
D41977 N41977 0 diode
R41978 N41977 N41978 10
D41978 N41978 0 diode
R41979 N41978 N41979 10
D41979 N41979 0 diode
R41980 N41979 N41980 10
D41980 N41980 0 diode
R41981 N41980 N41981 10
D41981 N41981 0 diode
R41982 N41981 N41982 10
D41982 N41982 0 diode
R41983 N41982 N41983 10
D41983 N41983 0 diode
R41984 N41983 N41984 10
D41984 N41984 0 diode
R41985 N41984 N41985 10
D41985 N41985 0 diode
R41986 N41985 N41986 10
D41986 N41986 0 diode
R41987 N41986 N41987 10
D41987 N41987 0 diode
R41988 N41987 N41988 10
D41988 N41988 0 diode
R41989 N41988 N41989 10
D41989 N41989 0 diode
R41990 N41989 N41990 10
D41990 N41990 0 diode
R41991 N41990 N41991 10
D41991 N41991 0 diode
R41992 N41991 N41992 10
D41992 N41992 0 diode
R41993 N41992 N41993 10
D41993 N41993 0 diode
R41994 N41993 N41994 10
D41994 N41994 0 diode
R41995 N41994 N41995 10
D41995 N41995 0 diode
R41996 N41995 N41996 10
D41996 N41996 0 diode
R41997 N41996 N41997 10
D41997 N41997 0 diode
R41998 N41997 N41998 10
D41998 N41998 0 diode
R41999 N41998 N41999 10
D41999 N41999 0 diode
R42000 N41999 N42000 10
D42000 N42000 0 diode
R42001 N42000 N42001 10
D42001 N42001 0 diode
R42002 N42001 N42002 10
D42002 N42002 0 diode
R42003 N42002 N42003 10
D42003 N42003 0 diode
R42004 N42003 N42004 10
D42004 N42004 0 diode
R42005 N42004 N42005 10
D42005 N42005 0 diode
R42006 N42005 N42006 10
D42006 N42006 0 diode
R42007 N42006 N42007 10
D42007 N42007 0 diode
R42008 N42007 N42008 10
D42008 N42008 0 diode
R42009 N42008 N42009 10
D42009 N42009 0 diode
R42010 N42009 N42010 10
D42010 N42010 0 diode
R42011 N42010 N42011 10
D42011 N42011 0 diode
R42012 N42011 N42012 10
D42012 N42012 0 diode
R42013 N42012 N42013 10
D42013 N42013 0 diode
R42014 N42013 N42014 10
D42014 N42014 0 diode
R42015 N42014 N42015 10
D42015 N42015 0 diode
R42016 N42015 N42016 10
D42016 N42016 0 diode
R42017 N42016 N42017 10
D42017 N42017 0 diode
R42018 N42017 N42018 10
D42018 N42018 0 diode
R42019 N42018 N42019 10
D42019 N42019 0 diode
R42020 N42019 N42020 10
D42020 N42020 0 diode
R42021 N42020 N42021 10
D42021 N42021 0 diode
R42022 N42021 N42022 10
D42022 N42022 0 diode
R42023 N42022 N42023 10
D42023 N42023 0 diode
R42024 N42023 N42024 10
D42024 N42024 0 diode
R42025 N42024 N42025 10
D42025 N42025 0 diode
R42026 N42025 N42026 10
D42026 N42026 0 diode
R42027 N42026 N42027 10
D42027 N42027 0 diode
R42028 N42027 N42028 10
D42028 N42028 0 diode
R42029 N42028 N42029 10
D42029 N42029 0 diode
R42030 N42029 N42030 10
D42030 N42030 0 diode
R42031 N42030 N42031 10
D42031 N42031 0 diode
R42032 N42031 N42032 10
D42032 N42032 0 diode
R42033 N42032 N42033 10
D42033 N42033 0 diode
R42034 N42033 N42034 10
D42034 N42034 0 diode
R42035 N42034 N42035 10
D42035 N42035 0 diode
R42036 N42035 N42036 10
D42036 N42036 0 diode
R42037 N42036 N42037 10
D42037 N42037 0 diode
R42038 N42037 N42038 10
D42038 N42038 0 diode
R42039 N42038 N42039 10
D42039 N42039 0 diode
R42040 N42039 N42040 10
D42040 N42040 0 diode
R42041 N42040 N42041 10
D42041 N42041 0 diode
R42042 N42041 N42042 10
D42042 N42042 0 diode
R42043 N42042 N42043 10
D42043 N42043 0 diode
R42044 N42043 N42044 10
D42044 N42044 0 diode
R42045 N42044 N42045 10
D42045 N42045 0 diode
R42046 N42045 N42046 10
D42046 N42046 0 diode
R42047 N42046 N42047 10
D42047 N42047 0 diode
R42048 N42047 N42048 10
D42048 N42048 0 diode
R42049 N42048 N42049 10
D42049 N42049 0 diode
R42050 N42049 N42050 10
D42050 N42050 0 diode
R42051 N42050 N42051 10
D42051 N42051 0 diode
R42052 N42051 N42052 10
D42052 N42052 0 diode
R42053 N42052 N42053 10
D42053 N42053 0 diode
R42054 N42053 N42054 10
D42054 N42054 0 diode
R42055 N42054 N42055 10
D42055 N42055 0 diode
R42056 N42055 N42056 10
D42056 N42056 0 diode
R42057 N42056 N42057 10
D42057 N42057 0 diode
R42058 N42057 N42058 10
D42058 N42058 0 diode
R42059 N42058 N42059 10
D42059 N42059 0 diode
R42060 N42059 N42060 10
D42060 N42060 0 diode
R42061 N42060 N42061 10
D42061 N42061 0 diode
R42062 N42061 N42062 10
D42062 N42062 0 diode
R42063 N42062 N42063 10
D42063 N42063 0 diode
R42064 N42063 N42064 10
D42064 N42064 0 diode
R42065 N42064 N42065 10
D42065 N42065 0 diode
R42066 N42065 N42066 10
D42066 N42066 0 diode
R42067 N42066 N42067 10
D42067 N42067 0 diode
R42068 N42067 N42068 10
D42068 N42068 0 diode
R42069 N42068 N42069 10
D42069 N42069 0 diode
R42070 N42069 N42070 10
D42070 N42070 0 diode
R42071 N42070 N42071 10
D42071 N42071 0 diode
R42072 N42071 N42072 10
D42072 N42072 0 diode
R42073 N42072 N42073 10
D42073 N42073 0 diode
R42074 N42073 N42074 10
D42074 N42074 0 diode
R42075 N42074 N42075 10
D42075 N42075 0 diode
R42076 N42075 N42076 10
D42076 N42076 0 diode
R42077 N42076 N42077 10
D42077 N42077 0 diode
R42078 N42077 N42078 10
D42078 N42078 0 diode
R42079 N42078 N42079 10
D42079 N42079 0 diode
R42080 N42079 N42080 10
D42080 N42080 0 diode
R42081 N42080 N42081 10
D42081 N42081 0 diode
R42082 N42081 N42082 10
D42082 N42082 0 diode
R42083 N42082 N42083 10
D42083 N42083 0 diode
R42084 N42083 N42084 10
D42084 N42084 0 diode
R42085 N42084 N42085 10
D42085 N42085 0 diode
R42086 N42085 N42086 10
D42086 N42086 0 diode
R42087 N42086 N42087 10
D42087 N42087 0 diode
R42088 N42087 N42088 10
D42088 N42088 0 diode
R42089 N42088 N42089 10
D42089 N42089 0 diode
R42090 N42089 N42090 10
D42090 N42090 0 diode
R42091 N42090 N42091 10
D42091 N42091 0 diode
R42092 N42091 N42092 10
D42092 N42092 0 diode
R42093 N42092 N42093 10
D42093 N42093 0 diode
R42094 N42093 N42094 10
D42094 N42094 0 diode
R42095 N42094 N42095 10
D42095 N42095 0 diode
R42096 N42095 N42096 10
D42096 N42096 0 diode
R42097 N42096 N42097 10
D42097 N42097 0 diode
R42098 N42097 N42098 10
D42098 N42098 0 diode
R42099 N42098 N42099 10
D42099 N42099 0 diode
R42100 N42099 N42100 10
D42100 N42100 0 diode
R42101 N42100 N42101 10
D42101 N42101 0 diode
R42102 N42101 N42102 10
D42102 N42102 0 diode
R42103 N42102 N42103 10
D42103 N42103 0 diode
R42104 N42103 N42104 10
D42104 N42104 0 diode
R42105 N42104 N42105 10
D42105 N42105 0 diode
R42106 N42105 N42106 10
D42106 N42106 0 diode
R42107 N42106 N42107 10
D42107 N42107 0 diode
R42108 N42107 N42108 10
D42108 N42108 0 diode
R42109 N42108 N42109 10
D42109 N42109 0 diode
R42110 N42109 N42110 10
D42110 N42110 0 diode
R42111 N42110 N42111 10
D42111 N42111 0 diode
R42112 N42111 N42112 10
D42112 N42112 0 diode
R42113 N42112 N42113 10
D42113 N42113 0 diode
R42114 N42113 N42114 10
D42114 N42114 0 diode
R42115 N42114 N42115 10
D42115 N42115 0 diode
R42116 N42115 N42116 10
D42116 N42116 0 diode
R42117 N42116 N42117 10
D42117 N42117 0 diode
R42118 N42117 N42118 10
D42118 N42118 0 diode
R42119 N42118 N42119 10
D42119 N42119 0 diode
R42120 N42119 N42120 10
D42120 N42120 0 diode
R42121 N42120 N42121 10
D42121 N42121 0 diode
R42122 N42121 N42122 10
D42122 N42122 0 diode
R42123 N42122 N42123 10
D42123 N42123 0 diode
R42124 N42123 N42124 10
D42124 N42124 0 diode
R42125 N42124 N42125 10
D42125 N42125 0 diode
R42126 N42125 N42126 10
D42126 N42126 0 diode
R42127 N42126 N42127 10
D42127 N42127 0 diode
R42128 N42127 N42128 10
D42128 N42128 0 diode
R42129 N42128 N42129 10
D42129 N42129 0 diode
R42130 N42129 N42130 10
D42130 N42130 0 diode
R42131 N42130 N42131 10
D42131 N42131 0 diode
R42132 N42131 N42132 10
D42132 N42132 0 diode
R42133 N42132 N42133 10
D42133 N42133 0 diode
R42134 N42133 N42134 10
D42134 N42134 0 diode
R42135 N42134 N42135 10
D42135 N42135 0 diode
R42136 N42135 N42136 10
D42136 N42136 0 diode
R42137 N42136 N42137 10
D42137 N42137 0 diode
R42138 N42137 N42138 10
D42138 N42138 0 diode
R42139 N42138 N42139 10
D42139 N42139 0 diode
R42140 N42139 N42140 10
D42140 N42140 0 diode
R42141 N42140 N42141 10
D42141 N42141 0 diode
R42142 N42141 N42142 10
D42142 N42142 0 diode
R42143 N42142 N42143 10
D42143 N42143 0 diode
R42144 N42143 N42144 10
D42144 N42144 0 diode
R42145 N42144 N42145 10
D42145 N42145 0 diode
R42146 N42145 N42146 10
D42146 N42146 0 diode
R42147 N42146 N42147 10
D42147 N42147 0 diode
R42148 N42147 N42148 10
D42148 N42148 0 diode
R42149 N42148 N42149 10
D42149 N42149 0 diode
R42150 N42149 N42150 10
D42150 N42150 0 diode
R42151 N42150 N42151 10
D42151 N42151 0 diode
R42152 N42151 N42152 10
D42152 N42152 0 diode
R42153 N42152 N42153 10
D42153 N42153 0 diode
R42154 N42153 N42154 10
D42154 N42154 0 diode
R42155 N42154 N42155 10
D42155 N42155 0 diode
R42156 N42155 N42156 10
D42156 N42156 0 diode
R42157 N42156 N42157 10
D42157 N42157 0 diode
R42158 N42157 N42158 10
D42158 N42158 0 diode
R42159 N42158 N42159 10
D42159 N42159 0 diode
R42160 N42159 N42160 10
D42160 N42160 0 diode
R42161 N42160 N42161 10
D42161 N42161 0 diode
R42162 N42161 N42162 10
D42162 N42162 0 diode
R42163 N42162 N42163 10
D42163 N42163 0 diode
R42164 N42163 N42164 10
D42164 N42164 0 diode
R42165 N42164 N42165 10
D42165 N42165 0 diode
R42166 N42165 N42166 10
D42166 N42166 0 diode
R42167 N42166 N42167 10
D42167 N42167 0 diode
R42168 N42167 N42168 10
D42168 N42168 0 diode
R42169 N42168 N42169 10
D42169 N42169 0 diode
R42170 N42169 N42170 10
D42170 N42170 0 diode
R42171 N42170 N42171 10
D42171 N42171 0 diode
R42172 N42171 N42172 10
D42172 N42172 0 diode
R42173 N42172 N42173 10
D42173 N42173 0 diode
R42174 N42173 N42174 10
D42174 N42174 0 diode
R42175 N42174 N42175 10
D42175 N42175 0 diode
R42176 N42175 N42176 10
D42176 N42176 0 diode
R42177 N42176 N42177 10
D42177 N42177 0 diode
R42178 N42177 N42178 10
D42178 N42178 0 diode
R42179 N42178 N42179 10
D42179 N42179 0 diode
R42180 N42179 N42180 10
D42180 N42180 0 diode
R42181 N42180 N42181 10
D42181 N42181 0 diode
R42182 N42181 N42182 10
D42182 N42182 0 diode
R42183 N42182 N42183 10
D42183 N42183 0 diode
R42184 N42183 N42184 10
D42184 N42184 0 diode
R42185 N42184 N42185 10
D42185 N42185 0 diode
R42186 N42185 N42186 10
D42186 N42186 0 diode
R42187 N42186 N42187 10
D42187 N42187 0 diode
R42188 N42187 N42188 10
D42188 N42188 0 diode
R42189 N42188 N42189 10
D42189 N42189 0 diode
R42190 N42189 N42190 10
D42190 N42190 0 diode
R42191 N42190 N42191 10
D42191 N42191 0 diode
R42192 N42191 N42192 10
D42192 N42192 0 diode
R42193 N42192 N42193 10
D42193 N42193 0 diode
R42194 N42193 N42194 10
D42194 N42194 0 diode
R42195 N42194 N42195 10
D42195 N42195 0 diode
R42196 N42195 N42196 10
D42196 N42196 0 diode
R42197 N42196 N42197 10
D42197 N42197 0 diode
R42198 N42197 N42198 10
D42198 N42198 0 diode
R42199 N42198 N42199 10
D42199 N42199 0 diode
R42200 N42199 N42200 10
D42200 N42200 0 diode
R42201 N42200 N42201 10
D42201 N42201 0 diode
R42202 N42201 N42202 10
D42202 N42202 0 diode
R42203 N42202 N42203 10
D42203 N42203 0 diode
R42204 N42203 N42204 10
D42204 N42204 0 diode
R42205 N42204 N42205 10
D42205 N42205 0 diode
R42206 N42205 N42206 10
D42206 N42206 0 diode
R42207 N42206 N42207 10
D42207 N42207 0 diode
R42208 N42207 N42208 10
D42208 N42208 0 diode
R42209 N42208 N42209 10
D42209 N42209 0 diode
R42210 N42209 N42210 10
D42210 N42210 0 diode
R42211 N42210 N42211 10
D42211 N42211 0 diode
R42212 N42211 N42212 10
D42212 N42212 0 diode
R42213 N42212 N42213 10
D42213 N42213 0 diode
R42214 N42213 N42214 10
D42214 N42214 0 diode
R42215 N42214 N42215 10
D42215 N42215 0 diode
R42216 N42215 N42216 10
D42216 N42216 0 diode
R42217 N42216 N42217 10
D42217 N42217 0 diode
R42218 N42217 N42218 10
D42218 N42218 0 diode
R42219 N42218 N42219 10
D42219 N42219 0 diode
R42220 N42219 N42220 10
D42220 N42220 0 diode
R42221 N42220 N42221 10
D42221 N42221 0 diode
R42222 N42221 N42222 10
D42222 N42222 0 diode
R42223 N42222 N42223 10
D42223 N42223 0 diode
R42224 N42223 N42224 10
D42224 N42224 0 diode
R42225 N42224 N42225 10
D42225 N42225 0 diode
R42226 N42225 N42226 10
D42226 N42226 0 diode
R42227 N42226 N42227 10
D42227 N42227 0 diode
R42228 N42227 N42228 10
D42228 N42228 0 diode
R42229 N42228 N42229 10
D42229 N42229 0 diode
R42230 N42229 N42230 10
D42230 N42230 0 diode
R42231 N42230 N42231 10
D42231 N42231 0 diode
R42232 N42231 N42232 10
D42232 N42232 0 diode
R42233 N42232 N42233 10
D42233 N42233 0 diode
R42234 N42233 N42234 10
D42234 N42234 0 diode
R42235 N42234 N42235 10
D42235 N42235 0 diode
R42236 N42235 N42236 10
D42236 N42236 0 diode
R42237 N42236 N42237 10
D42237 N42237 0 diode
R42238 N42237 N42238 10
D42238 N42238 0 diode
R42239 N42238 N42239 10
D42239 N42239 0 diode
R42240 N42239 N42240 10
D42240 N42240 0 diode
R42241 N42240 N42241 10
D42241 N42241 0 diode
R42242 N42241 N42242 10
D42242 N42242 0 diode
R42243 N42242 N42243 10
D42243 N42243 0 diode
R42244 N42243 N42244 10
D42244 N42244 0 diode
R42245 N42244 N42245 10
D42245 N42245 0 diode
R42246 N42245 N42246 10
D42246 N42246 0 diode
R42247 N42246 N42247 10
D42247 N42247 0 diode
R42248 N42247 N42248 10
D42248 N42248 0 diode
R42249 N42248 N42249 10
D42249 N42249 0 diode
R42250 N42249 N42250 10
D42250 N42250 0 diode
R42251 N42250 N42251 10
D42251 N42251 0 diode
R42252 N42251 N42252 10
D42252 N42252 0 diode
R42253 N42252 N42253 10
D42253 N42253 0 diode
R42254 N42253 N42254 10
D42254 N42254 0 diode
R42255 N42254 N42255 10
D42255 N42255 0 diode
R42256 N42255 N42256 10
D42256 N42256 0 diode
R42257 N42256 N42257 10
D42257 N42257 0 diode
R42258 N42257 N42258 10
D42258 N42258 0 diode
R42259 N42258 N42259 10
D42259 N42259 0 diode
R42260 N42259 N42260 10
D42260 N42260 0 diode
R42261 N42260 N42261 10
D42261 N42261 0 diode
R42262 N42261 N42262 10
D42262 N42262 0 diode
R42263 N42262 N42263 10
D42263 N42263 0 diode
R42264 N42263 N42264 10
D42264 N42264 0 diode
R42265 N42264 N42265 10
D42265 N42265 0 diode
R42266 N42265 N42266 10
D42266 N42266 0 diode
R42267 N42266 N42267 10
D42267 N42267 0 diode
R42268 N42267 N42268 10
D42268 N42268 0 diode
R42269 N42268 N42269 10
D42269 N42269 0 diode
R42270 N42269 N42270 10
D42270 N42270 0 diode
R42271 N42270 N42271 10
D42271 N42271 0 diode
R42272 N42271 N42272 10
D42272 N42272 0 diode
R42273 N42272 N42273 10
D42273 N42273 0 diode
R42274 N42273 N42274 10
D42274 N42274 0 diode
R42275 N42274 N42275 10
D42275 N42275 0 diode
R42276 N42275 N42276 10
D42276 N42276 0 diode
R42277 N42276 N42277 10
D42277 N42277 0 diode
R42278 N42277 N42278 10
D42278 N42278 0 diode
R42279 N42278 N42279 10
D42279 N42279 0 diode
R42280 N42279 N42280 10
D42280 N42280 0 diode
R42281 N42280 N42281 10
D42281 N42281 0 diode
R42282 N42281 N42282 10
D42282 N42282 0 diode
R42283 N42282 N42283 10
D42283 N42283 0 diode
R42284 N42283 N42284 10
D42284 N42284 0 diode
R42285 N42284 N42285 10
D42285 N42285 0 diode
R42286 N42285 N42286 10
D42286 N42286 0 diode
R42287 N42286 N42287 10
D42287 N42287 0 diode
R42288 N42287 N42288 10
D42288 N42288 0 diode
R42289 N42288 N42289 10
D42289 N42289 0 diode
R42290 N42289 N42290 10
D42290 N42290 0 diode
R42291 N42290 N42291 10
D42291 N42291 0 diode
R42292 N42291 N42292 10
D42292 N42292 0 diode
R42293 N42292 N42293 10
D42293 N42293 0 diode
R42294 N42293 N42294 10
D42294 N42294 0 diode
R42295 N42294 N42295 10
D42295 N42295 0 diode
R42296 N42295 N42296 10
D42296 N42296 0 diode
R42297 N42296 N42297 10
D42297 N42297 0 diode
R42298 N42297 N42298 10
D42298 N42298 0 diode
R42299 N42298 N42299 10
D42299 N42299 0 diode
R42300 N42299 N42300 10
D42300 N42300 0 diode
R42301 N42300 N42301 10
D42301 N42301 0 diode
R42302 N42301 N42302 10
D42302 N42302 0 diode
R42303 N42302 N42303 10
D42303 N42303 0 diode
R42304 N42303 N42304 10
D42304 N42304 0 diode
R42305 N42304 N42305 10
D42305 N42305 0 diode
R42306 N42305 N42306 10
D42306 N42306 0 diode
R42307 N42306 N42307 10
D42307 N42307 0 diode
R42308 N42307 N42308 10
D42308 N42308 0 diode
R42309 N42308 N42309 10
D42309 N42309 0 diode
R42310 N42309 N42310 10
D42310 N42310 0 diode
R42311 N42310 N42311 10
D42311 N42311 0 diode
R42312 N42311 N42312 10
D42312 N42312 0 diode
R42313 N42312 N42313 10
D42313 N42313 0 diode
R42314 N42313 N42314 10
D42314 N42314 0 diode
R42315 N42314 N42315 10
D42315 N42315 0 diode
R42316 N42315 N42316 10
D42316 N42316 0 diode
R42317 N42316 N42317 10
D42317 N42317 0 diode
R42318 N42317 N42318 10
D42318 N42318 0 diode
R42319 N42318 N42319 10
D42319 N42319 0 diode
R42320 N42319 N42320 10
D42320 N42320 0 diode
R42321 N42320 N42321 10
D42321 N42321 0 diode
R42322 N42321 N42322 10
D42322 N42322 0 diode
R42323 N42322 N42323 10
D42323 N42323 0 diode
R42324 N42323 N42324 10
D42324 N42324 0 diode
R42325 N42324 N42325 10
D42325 N42325 0 diode
R42326 N42325 N42326 10
D42326 N42326 0 diode
R42327 N42326 N42327 10
D42327 N42327 0 diode
R42328 N42327 N42328 10
D42328 N42328 0 diode
R42329 N42328 N42329 10
D42329 N42329 0 diode
R42330 N42329 N42330 10
D42330 N42330 0 diode
R42331 N42330 N42331 10
D42331 N42331 0 diode
R42332 N42331 N42332 10
D42332 N42332 0 diode
R42333 N42332 N42333 10
D42333 N42333 0 diode
R42334 N42333 N42334 10
D42334 N42334 0 diode
R42335 N42334 N42335 10
D42335 N42335 0 diode
R42336 N42335 N42336 10
D42336 N42336 0 diode
R42337 N42336 N42337 10
D42337 N42337 0 diode
R42338 N42337 N42338 10
D42338 N42338 0 diode
R42339 N42338 N42339 10
D42339 N42339 0 diode
R42340 N42339 N42340 10
D42340 N42340 0 diode
R42341 N42340 N42341 10
D42341 N42341 0 diode
R42342 N42341 N42342 10
D42342 N42342 0 diode
R42343 N42342 N42343 10
D42343 N42343 0 diode
R42344 N42343 N42344 10
D42344 N42344 0 diode
R42345 N42344 N42345 10
D42345 N42345 0 diode
R42346 N42345 N42346 10
D42346 N42346 0 diode
R42347 N42346 N42347 10
D42347 N42347 0 diode
R42348 N42347 N42348 10
D42348 N42348 0 diode
R42349 N42348 N42349 10
D42349 N42349 0 diode
R42350 N42349 N42350 10
D42350 N42350 0 diode
R42351 N42350 N42351 10
D42351 N42351 0 diode
R42352 N42351 N42352 10
D42352 N42352 0 diode
R42353 N42352 N42353 10
D42353 N42353 0 diode
R42354 N42353 N42354 10
D42354 N42354 0 diode
R42355 N42354 N42355 10
D42355 N42355 0 diode
R42356 N42355 N42356 10
D42356 N42356 0 diode
R42357 N42356 N42357 10
D42357 N42357 0 diode
R42358 N42357 N42358 10
D42358 N42358 0 diode
R42359 N42358 N42359 10
D42359 N42359 0 diode
R42360 N42359 N42360 10
D42360 N42360 0 diode
R42361 N42360 N42361 10
D42361 N42361 0 diode
R42362 N42361 N42362 10
D42362 N42362 0 diode
R42363 N42362 N42363 10
D42363 N42363 0 diode
R42364 N42363 N42364 10
D42364 N42364 0 diode
R42365 N42364 N42365 10
D42365 N42365 0 diode
R42366 N42365 N42366 10
D42366 N42366 0 diode
R42367 N42366 N42367 10
D42367 N42367 0 diode
R42368 N42367 N42368 10
D42368 N42368 0 diode
R42369 N42368 N42369 10
D42369 N42369 0 diode
R42370 N42369 N42370 10
D42370 N42370 0 diode
R42371 N42370 N42371 10
D42371 N42371 0 diode
R42372 N42371 N42372 10
D42372 N42372 0 diode
R42373 N42372 N42373 10
D42373 N42373 0 diode
R42374 N42373 N42374 10
D42374 N42374 0 diode
R42375 N42374 N42375 10
D42375 N42375 0 diode
R42376 N42375 N42376 10
D42376 N42376 0 diode
R42377 N42376 N42377 10
D42377 N42377 0 diode
R42378 N42377 N42378 10
D42378 N42378 0 diode
R42379 N42378 N42379 10
D42379 N42379 0 diode
R42380 N42379 N42380 10
D42380 N42380 0 diode
R42381 N42380 N42381 10
D42381 N42381 0 diode
R42382 N42381 N42382 10
D42382 N42382 0 diode
R42383 N42382 N42383 10
D42383 N42383 0 diode
R42384 N42383 N42384 10
D42384 N42384 0 diode
R42385 N42384 N42385 10
D42385 N42385 0 diode
R42386 N42385 N42386 10
D42386 N42386 0 diode
R42387 N42386 N42387 10
D42387 N42387 0 diode
R42388 N42387 N42388 10
D42388 N42388 0 diode
R42389 N42388 N42389 10
D42389 N42389 0 diode
R42390 N42389 N42390 10
D42390 N42390 0 diode
R42391 N42390 N42391 10
D42391 N42391 0 diode
R42392 N42391 N42392 10
D42392 N42392 0 diode
R42393 N42392 N42393 10
D42393 N42393 0 diode
R42394 N42393 N42394 10
D42394 N42394 0 diode
R42395 N42394 N42395 10
D42395 N42395 0 diode
R42396 N42395 N42396 10
D42396 N42396 0 diode
R42397 N42396 N42397 10
D42397 N42397 0 diode
R42398 N42397 N42398 10
D42398 N42398 0 diode
R42399 N42398 N42399 10
D42399 N42399 0 diode
R42400 N42399 N42400 10
D42400 N42400 0 diode
R42401 N42400 N42401 10
D42401 N42401 0 diode
R42402 N42401 N42402 10
D42402 N42402 0 diode
R42403 N42402 N42403 10
D42403 N42403 0 diode
R42404 N42403 N42404 10
D42404 N42404 0 diode
R42405 N42404 N42405 10
D42405 N42405 0 diode
R42406 N42405 N42406 10
D42406 N42406 0 diode
R42407 N42406 N42407 10
D42407 N42407 0 diode
R42408 N42407 N42408 10
D42408 N42408 0 diode
R42409 N42408 N42409 10
D42409 N42409 0 diode
R42410 N42409 N42410 10
D42410 N42410 0 diode
R42411 N42410 N42411 10
D42411 N42411 0 diode
R42412 N42411 N42412 10
D42412 N42412 0 diode
R42413 N42412 N42413 10
D42413 N42413 0 diode
R42414 N42413 N42414 10
D42414 N42414 0 diode
R42415 N42414 N42415 10
D42415 N42415 0 diode
R42416 N42415 N42416 10
D42416 N42416 0 diode
R42417 N42416 N42417 10
D42417 N42417 0 diode
R42418 N42417 N42418 10
D42418 N42418 0 diode
R42419 N42418 N42419 10
D42419 N42419 0 diode
R42420 N42419 N42420 10
D42420 N42420 0 diode
R42421 N42420 N42421 10
D42421 N42421 0 diode
R42422 N42421 N42422 10
D42422 N42422 0 diode
R42423 N42422 N42423 10
D42423 N42423 0 diode
R42424 N42423 N42424 10
D42424 N42424 0 diode
R42425 N42424 N42425 10
D42425 N42425 0 diode
R42426 N42425 N42426 10
D42426 N42426 0 diode
R42427 N42426 N42427 10
D42427 N42427 0 diode
R42428 N42427 N42428 10
D42428 N42428 0 diode
R42429 N42428 N42429 10
D42429 N42429 0 diode
R42430 N42429 N42430 10
D42430 N42430 0 diode
R42431 N42430 N42431 10
D42431 N42431 0 diode
R42432 N42431 N42432 10
D42432 N42432 0 diode
R42433 N42432 N42433 10
D42433 N42433 0 diode
R42434 N42433 N42434 10
D42434 N42434 0 diode
R42435 N42434 N42435 10
D42435 N42435 0 diode
R42436 N42435 N42436 10
D42436 N42436 0 diode
R42437 N42436 N42437 10
D42437 N42437 0 diode
R42438 N42437 N42438 10
D42438 N42438 0 diode
R42439 N42438 N42439 10
D42439 N42439 0 diode
R42440 N42439 N42440 10
D42440 N42440 0 diode
R42441 N42440 N42441 10
D42441 N42441 0 diode
R42442 N42441 N42442 10
D42442 N42442 0 diode
R42443 N42442 N42443 10
D42443 N42443 0 diode
R42444 N42443 N42444 10
D42444 N42444 0 diode
R42445 N42444 N42445 10
D42445 N42445 0 diode
R42446 N42445 N42446 10
D42446 N42446 0 diode
R42447 N42446 N42447 10
D42447 N42447 0 diode
R42448 N42447 N42448 10
D42448 N42448 0 diode
R42449 N42448 N42449 10
D42449 N42449 0 diode
R42450 N42449 N42450 10
D42450 N42450 0 diode
R42451 N42450 N42451 10
D42451 N42451 0 diode
R42452 N42451 N42452 10
D42452 N42452 0 diode
R42453 N42452 N42453 10
D42453 N42453 0 diode
R42454 N42453 N42454 10
D42454 N42454 0 diode
R42455 N42454 N42455 10
D42455 N42455 0 diode
R42456 N42455 N42456 10
D42456 N42456 0 diode
R42457 N42456 N42457 10
D42457 N42457 0 diode
R42458 N42457 N42458 10
D42458 N42458 0 diode
R42459 N42458 N42459 10
D42459 N42459 0 diode
R42460 N42459 N42460 10
D42460 N42460 0 diode
R42461 N42460 N42461 10
D42461 N42461 0 diode
R42462 N42461 N42462 10
D42462 N42462 0 diode
R42463 N42462 N42463 10
D42463 N42463 0 diode
R42464 N42463 N42464 10
D42464 N42464 0 diode
R42465 N42464 N42465 10
D42465 N42465 0 diode
R42466 N42465 N42466 10
D42466 N42466 0 diode
R42467 N42466 N42467 10
D42467 N42467 0 diode
R42468 N42467 N42468 10
D42468 N42468 0 diode
R42469 N42468 N42469 10
D42469 N42469 0 diode
R42470 N42469 N42470 10
D42470 N42470 0 diode
R42471 N42470 N42471 10
D42471 N42471 0 diode
R42472 N42471 N42472 10
D42472 N42472 0 diode
R42473 N42472 N42473 10
D42473 N42473 0 diode
R42474 N42473 N42474 10
D42474 N42474 0 diode
R42475 N42474 N42475 10
D42475 N42475 0 diode
R42476 N42475 N42476 10
D42476 N42476 0 diode
R42477 N42476 N42477 10
D42477 N42477 0 diode
R42478 N42477 N42478 10
D42478 N42478 0 diode
R42479 N42478 N42479 10
D42479 N42479 0 diode
R42480 N42479 N42480 10
D42480 N42480 0 diode
R42481 N42480 N42481 10
D42481 N42481 0 diode
R42482 N42481 N42482 10
D42482 N42482 0 diode
R42483 N42482 N42483 10
D42483 N42483 0 diode
R42484 N42483 N42484 10
D42484 N42484 0 diode
R42485 N42484 N42485 10
D42485 N42485 0 diode
R42486 N42485 N42486 10
D42486 N42486 0 diode
R42487 N42486 N42487 10
D42487 N42487 0 diode
R42488 N42487 N42488 10
D42488 N42488 0 diode
R42489 N42488 N42489 10
D42489 N42489 0 diode
R42490 N42489 N42490 10
D42490 N42490 0 diode
R42491 N42490 N42491 10
D42491 N42491 0 diode
R42492 N42491 N42492 10
D42492 N42492 0 diode
R42493 N42492 N42493 10
D42493 N42493 0 diode
R42494 N42493 N42494 10
D42494 N42494 0 diode
R42495 N42494 N42495 10
D42495 N42495 0 diode
R42496 N42495 N42496 10
D42496 N42496 0 diode
R42497 N42496 N42497 10
D42497 N42497 0 diode
R42498 N42497 N42498 10
D42498 N42498 0 diode
R42499 N42498 N42499 10
D42499 N42499 0 diode
R42500 N42499 N42500 10
D42500 N42500 0 diode
R42501 N42500 N42501 10
D42501 N42501 0 diode
R42502 N42501 N42502 10
D42502 N42502 0 diode
R42503 N42502 N42503 10
D42503 N42503 0 diode
R42504 N42503 N42504 10
D42504 N42504 0 diode
R42505 N42504 N42505 10
D42505 N42505 0 diode
R42506 N42505 N42506 10
D42506 N42506 0 diode
R42507 N42506 N42507 10
D42507 N42507 0 diode
R42508 N42507 N42508 10
D42508 N42508 0 diode
R42509 N42508 N42509 10
D42509 N42509 0 diode
R42510 N42509 N42510 10
D42510 N42510 0 diode
R42511 N42510 N42511 10
D42511 N42511 0 diode
R42512 N42511 N42512 10
D42512 N42512 0 diode
R42513 N42512 N42513 10
D42513 N42513 0 diode
R42514 N42513 N42514 10
D42514 N42514 0 diode
R42515 N42514 N42515 10
D42515 N42515 0 diode
R42516 N42515 N42516 10
D42516 N42516 0 diode
R42517 N42516 N42517 10
D42517 N42517 0 diode
R42518 N42517 N42518 10
D42518 N42518 0 diode
R42519 N42518 N42519 10
D42519 N42519 0 diode
R42520 N42519 N42520 10
D42520 N42520 0 diode
R42521 N42520 N42521 10
D42521 N42521 0 diode
R42522 N42521 N42522 10
D42522 N42522 0 diode
R42523 N42522 N42523 10
D42523 N42523 0 diode
R42524 N42523 N42524 10
D42524 N42524 0 diode
R42525 N42524 N42525 10
D42525 N42525 0 diode
R42526 N42525 N42526 10
D42526 N42526 0 diode
R42527 N42526 N42527 10
D42527 N42527 0 diode
R42528 N42527 N42528 10
D42528 N42528 0 diode
R42529 N42528 N42529 10
D42529 N42529 0 diode
R42530 N42529 N42530 10
D42530 N42530 0 diode
R42531 N42530 N42531 10
D42531 N42531 0 diode
R42532 N42531 N42532 10
D42532 N42532 0 diode
R42533 N42532 N42533 10
D42533 N42533 0 diode
R42534 N42533 N42534 10
D42534 N42534 0 diode
R42535 N42534 N42535 10
D42535 N42535 0 diode
R42536 N42535 N42536 10
D42536 N42536 0 diode
R42537 N42536 N42537 10
D42537 N42537 0 diode
R42538 N42537 N42538 10
D42538 N42538 0 diode
R42539 N42538 N42539 10
D42539 N42539 0 diode
R42540 N42539 N42540 10
D42540 N42540 0 diode
R42541 N42540 N42541 10
D42541 N42541 0 diode
R42542 N42541 N42542 10
D42542 N42542 0 diode
R42543 N42542 N42543 10
D42543 N42543 0 diode
R42544 N42543 N42544 10
D42544 N42544 0 diode
R42545 N42544 N42545 10
D42545 N42545 0 diode
R42546 N42545 N42546 10
D42546 N42546 0 diode
R42547 N42546 N42547 10
D42547 N42547 0 diode
R42548 N42547 N42548 10
D42548 N42548 0 diode
R42549 N42548 N42549 10
D42549 N42549 0 diode
R42550 N42549 N42550 10
D42550 N42550 0 diode
R42551 N42550 N42551 10
D42551 N42551 0 diode
R42552 N42551 N42552 10
D42552 N42552 0 diode
R42553 N42552 N42553 10
D42553 N42553 0 diode
R42554 N42553 N42554 10
D42554 N42554 0 diode
R42555 N42554 N42555 10
D42555 N42555 0 diode
R42556 N42555 N42556 10
D42556 N42556 0 diode
R42557 N42556 N42557 10
D42557 N42557 0 diode
R42558 N42557 N42558 10
D42558 N42558 0 diode
R42559 N42558 N42559 10
D42559 N42559 0 diode
R42560 N42559 N42560 10
D42560 N42560 0 diode
R42561 N42560 N42561 10
D42561 N42561 0 diode
R42562 N42561 N42562 10
D42562 N42562 0 diode
R42563 N42562 N42563 10
D42563 N42563 0 diode
R42564 N42563 N42564 10
D42564 N42564 0 diode
R42565 N42564 N42565 10
D42565 N42565 0 diode
R42566 N42565 N42566 10
D42566 N42566 0 diode
R42567 N42566 N42567 10
D42567 N42567 0 diode
R42568 N42567 N42568 10
D42568 N42568 0 diode
R42569 N42568 N42569 10
D42569 N42569 0 diode
R42570 N42569 N42570 10
D42570 N42570 0 diode
R42571 N42570 N42571 10
D42571 N42571 0 diode
R42572 N42571 N42572 10
D42572 N42572 0 diode
R42573 N42572 N42573 10
D42573 N42573 0 diode
R42574 N42573 N42574 10
D42574 N42574 0 diode
R42575 N42574 N42575 10
D42575 N42575 0 diode
R42576 N42575 N42576 10
D42576 N42576 0 diode
R42577 N42576 N42577 10
D42577 N42577 0 diode
R42578 N42577 N42578 10
D42578 N42578 0 diode
R42579 N42578 N42579 10
D42579 N42579 0 diode
R42580 N42579 N42580 10
D42580 N42580 0 diode
R42581 N42580 N42581 10
D42581 N42581 0 diode
R42582 N42581 N42582 10
D42582 N42582 0 diode
R42583 N42582 N42583 10
D42583 N42583 0 diode
R42584 N42583 N42584 10
D42584 N42584 0 diode
R42585 N42584 N42585 10
D42585 N42585 0 diode
R42586 N42585 N42586 10
D42586 N42586 0 diode
R42587 N42586 N42587 10
D42587 N42587 0 diode
R42588 N42587 N42588 10
D42588 N42588 0 diode
R42589 N42588 N42589 10
D42589 N42589 0 diode
R42590 N42589 N42590 10
D42590 N42590 0 diode
R42591 N42590 N42591 10
D42591 N42591 0 diode
R42592 N42591 N42592 10
D42592 N42592 0 diode
R42593 N42592 N42593 10
D42593 N42593 0 diode
R42594 N42593 N42594 10
D42594 N42594 0 diode
R42595 N42594 N42595 10
D42595 N42595 0 diode
R42596 N42595 N42596 10
D42596 N42596 0 diode
R42597 N42596 N42597 10
D42597 N42597 0 diode
R42598 N42597 N42598 10
D42598 N42598 0 diode
R42599 N42598 N42599 10
D42599 N42599 0 diode
R42600 N42599 N42600 10
D42600 N42600 0 diode
R42601 N42600 N42601 10
D42601 N42601 0 diode
R42602 N42601 N42602 10
D42602 N42602 0 diode
R42603 N42602 N42603 10
D42603 N42603 0 diode
R42604 N42603 N42604 10
D42604 N42604 0 diode
R42605 N42604 N42605 10
D42605 N42605 0 diode
R42606 N42605 N42606 10
D42606 N42606 0 diode
R42607 N42606 N42607 10
D42607 N42607 0 diode
R42608 N42607 N42608 10
D42608 N42608 0 diode
R42609 N42608 N42609 10
D42609 N42609 0 diode
R42610 N42609 N42610 10
D42610 N42610 0 diode
R42611 N42610 N42611 10
D42611 N42611 0 diode
R42612 N42611 N42612 10
D42612 N42612 0 diode
R42613 N42612 N42613 10
D42613 N42613 0 diode
R42614 N42613 N42614 10
D42614 N42614 0 diode
R42615 N42614 N42615 10
D42615 N42615 0 diode
R42616 N42615 N42616 10
D42616 N42616 0 diode
R42617 N42616 N42617 10
D42617 N42617 0 diode
R42618 N42617 N42618 10
D42618 N42618 0 diode
R42619 N42618 N42619 10
D42619 N42619 0 diode
R42620 N42619 N42620 10
D42620 N42620 0 diode
R42621 N42620 N42621 10
D42621 N42621 0 diode
R42622 N42621 N42622 10
D42622 N42622 0 diode
R42623 N42622 N42623 10
D42623 N42623 0 diode
R42624 N42623 N42624 10
D42624 N42624 0 diode
R42625 N42624 N42625 10
D42625 N42625 0 diode
R42626 N42625 N42626 10
D42626 N42626 0 diode
R42627 N42626 N42627 10
D42627 N42627 0 diode
R42628 N42627 N42628 10
D42628 N42628 0 diode
R42629 N42628 N42629 10
D42629 N42629 0 diode
R42630 N42629 N42630 10
D42630 N42630 0 diode
R42631 N42630 N42631 10
D42631 N42631 0 diode
R42632 N42631 N42632 10
D42632 N42632 0 diode
R42633 N42632 N42633 10
D42633 N42633 0 diode
R42634 N42633 N42634 10
D42634 N42634 0 diode
R42635 N42634 N42635 10
D42635 N42635 0 diode
R42636 N42635 N42636 10
D42636 N42636 0 diode
R42637 N42636 N42637 10
D42637 N42637 0 diode
R42638 N42637 N42638 10
D42638 N42638 0 diode
R42639 N42638 N42639 10
D42639 N42639 0 diode
R42640 N42639 N42640 10
D42640 N42640 0 diode
R42641 N42640 N42641 10
D42641 N42641 0 diode
R42642 N42641 N42642 10
D42642 N42642 0 diode
R42643 N42642 N42643 10
D42643 N42643 0 diode
R42644 N42643 N42644 10
D42644 N42644 0 diode
R42645 N42644 N42645 10
D42645 N42645 0 diode
R42646 N42645 N42646 10
D42646 N42646 0 diode
R42647 N42646 N42647 10
D42647 N42647 0 diode
R42648 N42647 N42648 10
D42648 N42648 0 diode
R42649 N42648 N42649 10
D42649 N42649 0 diode
R42650 N42649 N42650 10
D42650 N42650 0 diode
R42651 N42650 N42651 10
D42651 N42651 0 diode
R42652 N42651 N42652 10
D42652 N42652 0 diode
R42653 N42652 N42653 10
D42653 N42653 0 diode
R42654 N42653 N42654 10
D42654 N42654 0 diode
R42655 N42654 N42655 10
D42655 N42655 0 diode
R42656 N42655 N42656 10
D42656 N42656 0 diode
R42657 N42656 N42657 10
D42657 N42657 0 diode
R42658 N42657 N42658 10
D42658 N42658 0 diode
R42659 N42658 N42659 10
D42659 N42659 0 diode
R42660 N42659 N42660 10
D42660 N42660 0 diode
R42661 N42660 N42661 10
D42661 N42661 0 diode
R42662 N42661 N42662 10
D42662 N42662 0 diode
R42663 N42662 N42663 10
D42663 N42663 0 diode
R42664 N42663 N42664 10
D42664 N42664 0 diode
R42665 N42664 N42665 10
D42665 N42665 0 diode
R42666 N42665 N42666 10
D42666 N42666 0 diode
R42667 N42666 N42667 10
D42667 N42667 0 diode
R42668 N42667 N42668 10
D42668 N42668 0 diode
R42669 N42668 N42669 10
D42669 N42669 0 diode
R42670 N42669 N42670 10
D42670 N42670 0 diode
R42671 N42670 N42671 10
D42671 N42671 0 diode
R42672 N42671 N42672 10
D42672 N42672 0 diode
R42673 N42672 N42673 10
D42673 N42673 0 diode
R42674 N42673 N42674 10
D42674 N42674 0 diode
R42675 N42674 N42675 10
D42675 N42675 0 diode
R42676 N42675 N42676 10
D42676 N42676 0 diode
R42677 N42676 N42677 10
D42677 N42677 0 diode
R42678 N42677 N42678 10
D42678 N42678 0 diode
R42679 N42678 N42679 10
D42679 N42679 0 diode
R42680 N42679 N42680 10
D42680 N42680 0 diode
R42681 N42680 N42681 10
D42681 N42681 0 diode
R42682 N42681 N42682 10
D42682 N42682 0 diode
R42683 N42682 N42683 10
D42683 N42683 0 diode
R42684 N42683 N42684 10
D42684 N42684 0 diode
R42685 N42684 N42685 10
D42685 N42685 0 diode
R42686 N42685 N42686 10
D42686 N42686 0 diode
R42687 N42686 N42687 10
D42687 N42687 0 diode
R42688 N42687 N42688 10
D42688 N42688 0 diode
R42689 N42688 N42689 10
D42689 N42689 0 diode
R42690 N42689 N42690 10
D42690 N42690 0 diode
R42691 N42690 N42691 10
D42691 N42691 0 diode
R42692 N42691 N42692 10
D42692 N42692 0 diode
R42693 N42692 N42693 10
D42693 N42693 0 diode
R42694 N42693 N42694 10
D42694 N42694 0 diode
R42695 N42694 N42695 10
D42695 N42695 0 diode
R42696 N42695 N42696 10
D42696 N42696 0 diode
R42697 N42696 N42697 10
D42697 N42697 0 diode
R42698 N42697 N42698 10
D42698 N42698 0 diode
R42699 N42698 N42699 10
D42699 N42699 0 diode
R42700 N42699 N42700 10
D42700 N42700 0 diode
R42701 N42700 N42701 10
D42701 N42701 0 diode
R42702 N42701 N42702 10
D42702 N42702 0 diode
R42703 N42702 N42703 10
D42703 N42703 0 diode
R42704 N42703 N42704 10
D42704 N42704 0 diode
R42705 N42704 N42705 10
D42705 N42705 0 diode
R42706 N42705 N42706 10
D42706 N42706 0 diode
R42707 N42706 N42707 10
D42707 N42707 0 diode
R42708 N42707 N42708 10
D42708 N42708 0 diode
R42709 N42708 N42709 10
D42709 N42709 0 diode
R42710 N42709 N42710 10
D42710 N42710 0 diode
R42711 N42710 N42711 10
D42711 N42711 0 diode
R42712 N42711 N42712 10
D42712 N42712 0 diode
R42713 N42712 N42713 10
D42713 N42713 0 diode
R42714 N42713 N42714 10
D42714 N42714 0 diode
R42715 N42714 N42715 10
D42715 N42715 0 diode
R42716 N42715 N42716 10
D42716 N42716 0 diode
R42717 N42716 N42717 10
D42717 N42717 0 diode
R42718 N42717 N42718 10
D42718 N42718 0 diode
R42719 N42718 N42719 10
D42719 N42719 0 diode
R42720 N42719 N42720 10
D42720 N42720 0 diode
R42721 N42720 N42721 10
D42721 N42721 0 diode
R42722 N42721 N42722 10
D42722 N42722 0 diode
R42723 N42722 N42723 10
D42723 N42723 0 diode
R42724 N42723 N42724 10
D42724 N42724 0 diode
R42725 N42724 N42725 10
D42725 N42725 0 diode
R42726 N42725 N42726 10
D42726 N42726 0 diode
R42727 N42726 N42727 10
D42727 N42727 0 diode
R42728 N42727 N42728 10
D42728 N42728 0 diode
R42729 N42728 N42729 10
D42729 N42729 0 diode
R42730 N42729 N42730 10
D42730 N42730 0 diode
R42731 N42730 N42731 10
D42731 N42731 0 diode
R42732 N42731 N42732 10
D42732 N42732 0 diode
R42733 N42732 N42733 10
D42733 N42733 0 diode
R42734 N42733 N42734 10
D42734 N42734 0 diode
R42735 N42734 N42735 10
D42735 N42735 0 diode
R42736 N42735 N42736 10
D42736 N42736 0 diode
R42737 N42736 N42737 10
D42737 N42737 0 diode
R42738 N42737 N42738 10
D42738 N42738 0 diode
R42739 N42738 N42739 10
D42739 N42739 0 diode
R42740 N42739 N42740 10
D42740 N42740 0 diode
R42741 N42740 N42741 10
D42741 N42741 0 diode
R42742 N42741 N42742 10
D42742 N42742 0 diode
R42743 N42742 N42743 10
D42743 N42743 0 diode
R42744 N42743 N42744 10
D42744 N42744 0 diode
R42745 N42744 N42745 10
D42745 N42745 0 diode
R42746 N42745 N42746 10
D42746 N42746 0 diode
R42747 N42746 N42747 10
D42747 N42747 0 diode
R42748 N42747 N42748 10
D42748 N42748 0 diode
R42749 N42748 N42749 10
D42749 N42749 0 diode
R42750 N42749 N42750 10
D42750 N42750 0 diode
R42751 N42750 N42751 10
D42751 N42751 0 diode
R42752 N42751 N42752 10
D42752 N42752 0 diode
R42753 N42752 N42753 10
D42753 N42753 0 diode
R42754 N42753 N42754 10
D42754 N42754 0 diode
R42755 N42754 N42755 10
D42755 N42755 0 diode
R42756 N42755 N42756 10
D42756 N42756 0 diode
R42757 N42756 N42757 10
D42757 N42757 0 diode
R42758 N42757 N42758 10
D42758 N42758 0 diode
R42759 N42758 N42759 10
D42759 N42759 0 diode
R42760 N42759 N42760 10
D42760 N42760 0 diode
R42761 N42760 N42761 10
D42761 N42761 0 diode
R42762 N42761 N42762 10
D42762 N42762 0 diode
R42763 N42762 N42763 10
D42763 N42763 0 diode
R42764 N42763 N42764 10
D42764 N42764 0 diode
R42765 N42764 N42765 10
D42765 N42765 0 diode
R42766 N42765 N42766 10
D42766 N42766 0 diode
R42767 N42766 N42767 10
D42767 N42767 0 diode
R42768 N42767 N42768 10
D42768 N42768 0 diode
R42769 N42768 N42769 10
D42769 N42769 0 diode
R42770 N42769 N42770 10
D42770 N42770 0 diode
R42771 N42770 N42771 10
D42771 N42771 0 diode
R42772 N42771 N42772 10
D42772 N42772 0 diode
R42773 N42772 N42773 10
D42773 N42773 0 diode
R42774 N42773 N42774 10
D42774 N42774 0 diode
R42775 N42774 N42775 10
D42775 N42775 0 diode
R42776 N42775 N42776 10
D42776 N42776 0 diode
R42777 N42776 N42777 10
D42777 N42777 0 diode
R42778 N42777 N42778 10
D42778 N42778 0 diode
R42779 N42778 N42779 10
D42779 N42779 0 diode
R42780 N42779 N42780 10
D42780 N42780 0 diode
R42781 N42780 N42781 10
D42781 N42781 0 diode
R42782 N42781 N42782 10
D42782 N42782 0 diode
R42783 N42782 N42783 10
D42783 N42783 0 diode
R42784 N42783 N42784 10
D42784 N42784 0 diode
R42785 N42784 N42785 10
D42785 N42785 0 diode
R42786 N42785 N42786 10
D42786 N42786 0 diode
R42787 N42786 N42787 10
D42787 N42787 0 diode
R42788 N42787 N42788 10
D42788 N42788 0 diode
R42789 N42788 N42789 10
D42789 N42789 0 diode
R42790 N42789 N42790 10
D42790 N42790 0 diode
R42791 N42790 N42791 10
D42791 N42791 0 diode
R42792 N42791 N42792 10
D42792 N42792 0 diode
R42793 N42792 N42793 10
D42793 N42793 0 diode
R42794 N42793 N42794 10
D42794 N42794 0 diode
R42795 N42794 N42795 10
D42795 N42795 0 diode
R42796 N42795 N42796 10
D42796 N42796 0 diode
R42797 N42796 N42797 10
D42797 N42797 0 diode
R42798 N42797 N42798 10
D42798 N42798 0 diode
R42799 N42798 N42799 10
D42799 N42799 0 diode
R42800 N42799 N42800 10
D42800 N42800 0 diode
R42801 N42800 N42801 10
D42801 N42801 0 diode
R42802 N42801 N42802 10
D42802 N42802 0 diode
R42803 N42802 N42803 10
D42803 N42803 0 diode
R42804 N42803 N42804 10
D42804 N42804 0 diode
R42805 N42804 N42805 10
D42805 N42805 0 diode
R42806 N42805 N42806 10
D42806 N42806 0 diode
R42807 N42806 N42807 10
D42807 N42807 0 diode
R42808 N42807 N42808 10
D42808 N42808 0 diode
R42809 N42808 N42809 10
D42809 N42809 0 diode
R42810 N42809 N42810 10
D42810 N42810 0 diode
R42811 N42810 N42811 10
D42811 N42811 0 diode
R42812 N42811 N42812 10
D42812 N42812 0 diode
R42813 N42812 N42813 10
D42813 N42813 0 diode
R42814 N42813 N42814 10
D42814 N42814 0 diode
R42815 N42814 N42815 10
D42815 N42815 0 diode
R42816 N42815 N42816 10
D42816 N42816 0 diode
R42817 N42816 N42817 10
D42817 N42817 0 diode
R42818 N42817 N42818 10
D42818 N42818 0 diode
R42819 N42818 N42819 10
D42819 N42819 0 diode
R42820 N42819 N42820 10
D42820 N42820 0 diode
R42821 N42820 N42821 10
D42821 N42821 0 diode
R42822 N42821 N42822 10
D42822 N42822 0 diode
R42823 N42822 N42823 10
D42823 N42823 0 diode
R42824 N42823 N42824 10
D42824 N42824 0 diode
R42825 N42824 N42825 10
D42825 N42825 0 diode
R42826 N42825 N42826 10
D42826 N42826 0 diode
R42827 N42826 N42827 10
D42827 N42827 0 diode
R42828 N42827 N42828 10
D42828 N42828 0 diode
R42829 N42828 N42829 10
D42829 N42829 0 diode
R42830 N42829 N42830 10
D42830 N42830 0 diode
R42831 N42830 N42831 10
D42831 N42831 0 diode
R42832 N42831 N42832 10
D42832 N42832 0 diode
R42833 N42832 N42833 10
D42833 N42833 0 diode
R42834 N42833 N42834 10
D42834 N42834 0 diode
R42835 N42834 N42835 10
D42835 N42835 0 diode
R42836 N42835 N42836 10
D42836 N42836 0 diode
R42837 N42836 N42837 10
D42837 N42837 0 diode
R42838 N42837 N42838 10
D42838 N42838 0 diode
R42839 N42838 N42839 10
D42839 N42839 0 diode
R42840 N42839 N42840 10
D42840 N42840 0 diode
R42841 N42840 N42841 10
D42841 N42841 0 diode
R42842 N42841 N42842 10
D42842 N42842 0 diode
R42843 N42842 N42843 10
D42843 N42843 0 diode
R42844 N42843 N42844 10
D42844 N42844 0 diode
R42845 N42844 N42845 10
D42845 N42845 0 diode
R42846 N42845 N42846 10
D42846 N42846 0 diode
R42847 N42846 N42847 10
D42847 N42847 0 diode
R42848 N42847 N42848 10
D42848 N42848 0 diode
R42849 N42848 N42849 10
D42849 N42849 0 diode
R42850 N42849 N42850 10
D42850 N42850 0 diode
R42851 N42850 N42851 10
D42851 N42851 0 diode
R42852 N42851 N42852 10
D42852 N42852 0 diode
R42853 N42852 N42853 10
D42853 N42853 0 diode
R42854 N42853 N42854 10
D42854 N42854 0 diode
R42855 N42854 N42855 10
D42855 N42855 0 diode
R42856 N42855 N42856 10
D42856 N42856 0 diode
R42857 N42856 N42857 10
D42857 N42857 0 diode
R42858 N42857 N42858 10
D42858 N42858 0 diode
R42859 N42858 N42859 10
D42859 N42859 0 diode
R42860 N42859 N42860 10
D42860 N42860 0 diode
R42861 N42860 N42861 10
D42861 N42861 0 diode
R42862 N42861 N42862 10
D42862 N42862 0 diode
R42863 N42862 N42863 10
D42863 N42863 0 diode
R42864 N42863 N42864 10
D42864 N42864 0 diode
R42865 N42864 N42865 10
D42865 N42865 0 diode
R42866 N42865 N42866 10
D42866 N42866 0 diode
R42867 N42866 N42867 10
D42867 N42867 0 diode
R42868 N42867 N42868 10
D42868 N42868 0 diode
R42869 N42868 N42869 10
D42869 N42869 0 diode
R42870 N42869 N42870 10
D42870 N42870 0 diode
R42871 N42870 N42871 10
D42871 N42871 0 diode
R42872 N42871 N42872 10
D42872 N42872 0 diode
R42873 N42872 N42873 10
D42873 N42873 0 diode
R42874 N42873 N42874 10
D42874 N42874 0 diode
R42875 N42874 N42875 10
D42875 N42875 0 diode
R42876 N42875 N42876 10
D42876 N42876 0 diode
R42877 N42876 N42877 10
D42877 N42877 0 diode
R42878 N42877 N42878 10
D42878 N42878 0 diode
R42879 N42878 N42879 10
D42879 N42879 0 diode
R42880 N42879 N42880 10
D42880 N42880 0 diode
R42881 N42880 N42881 10
D42881 N42881 0 diode
R42882 N42881 N42882 10
D42882 N42882 0 diode
R42883 N42882 N42883 10
D42883 N42883 0 diode
R42884 N42883 N42884 10
D42884 N42884 0 diode
R42885 N42884 N42885 10
D42885 N42885 0 diode
R42886 N42885 N42886 10
D42886 N42886 0 diode
R42887 N42886 N42887 10
D42887 N42887 0 diode
R42888 N42887 N42888 10
D42888 N42888 0 diode
R42889 N42888 N42889 10
D42889 N42889 0 diode
R42890 N42889 N42890 10
D42890 N42890 0 diode
R42891 N42890 N42891 10
D42891 N42891 0 diode
R42892 N42891 N42892 10
D42892 N42892 0 diode
R42893 N42892 N42893 10
D42893 N42893 0 diode
R42894 N42893 N42894 10
D42894 N42894 0 diode
R42895 N42894 N42895 10
D42895 N42895 0 diode
R42896 N42895 N42896 10
D42896 N42896 0 diode
R42897 N42896 N42897 10
D42897 N42897 0 diode
R42898 N42897 N42898 10
D42898 N42898 0 diode
R42899 N42898 N42899 10
D42899 N42899 0 diode
R42900 N42899 N42900 10
D42900 N42900 0 diode
R42901 N42900 N42901 10
D42901 N42901 0 diode
R42902 N42901 N42902 10
D42902 N42902 0 diode
R42903 N42902 N42903 10
D42903 N42903 0 diode
R42904 N42903 N42904 10
D42904 N42904 0 diode
R42905 N42904 N42905 10
D42905 N42905 0 diode
R42906 N42905 N42906 10
D42906 N42906 0 diode
R42907 N42906 N42907 10
D42907 N42907 0 diode
R42908 N42907 N42908 10
D42908 N42908 0 diode
R42909 N42908 N42909 10
D42909 N42909 0 diode
R42910 N42909 N42910 10
D42910 N42910 0 diode
R42911 N42910 N42911 10
D42911 N42911 0 diode
R42912 N42911 N42912 10
D42912 N42912 0 diode
R42913 N42912 N42913 10
D42913 N42913 0 diode
R42914 N42913 N42914 10
D42914 N42914 0 diode
R42915 N42914 N42915 10
D42915 N42915 0 diode
R42916 N42915 N42916 10
D42916 N42916 0 diode
R42917 N42916 N42917 10
D42917 N42917 0 diode
R42918 N42917 N42918 10
D42918 N42918 0 diode
R42919 N42918 N42919 10
D42919 N42919 0 diode
R42920 N42919 N42920 10
D42920 N42920 0 diode
R42921 N42920 N42921 10
D42921 N42921 0 diode
R42922 N42921 N42922 10
D42922 N42922 0 diode
R42923 N42922 N42923 10
D42923 N42923 0 diode
R42924 N42923 N42924 10
D42924 N42924 0 diode
R42925 N42924 N42925 10
D42925 N42925 0 diode
R42926 N42925 N42926 10
D42926 N42926 0 diode
R42927 N42926 N42927 10
D42927 N42927 0 diode
R42928 N42927 N42928 10
D42928 N42928 0 diode
R42929 N42928 N42929 10
D42929 N42929 0 diode
R42930 N42929 N42930 10
D42930 N42930 0 diode
R42931 N42930 N42931 10
D42931 N42931 0 diode
R42932 N42931 N42932 10
D42932 N42932 0 diode
R42933 N42932 N42933 10
D42933 N42933 0 diode
R42934 N42933 N42934 10
D42934 N42934 0 diode
R42935 N42934 N42935 10
D42935 N42935 0 diode
R42936 N42935 N42936 10
D42936 N42936 0 diode
R42937 N42936 N42937 10
D42937 N42937 0 diode
R42938 N42937 N42938 10
D42938 N42938 0 diode
R42939 N42938 N42939 10
D42939 N42939 0 diode
R42940 N42939 N42940 10
D42940 N42940 0 diode
R42941 N42940 N42941 10
D42941 N42941 0 diode
R42942 N42941 N42942 10
D42942 N42942 0 diode
R42943 N42942 N42943 10
D42943 N42943 0 diode
R42944 N42943 N42944 10
D42944 N42944 0 diode
R42945 N42944 N42945 10
D42945 N42945 0 diode
R42946 N42945 N42946 10
D42946 N42946 0 diode
R42947 N42946 N42947 10
D42947 N42947 0 diode
R42948 N42947 N42948 10
D42948 N42948 0 diode
R42949 N42948 N42949 10
D42949 N42949 0 diode
R42950 N42949 N42950 10
D42950 N42950 0 diode
R42951 N42950 N42951 10
D42951 N42951 0 diode
R42952 N42951 N42952 10
D42952 N42952 0 diode
R42953 N42952 N42953 10
D42953 N42953 0 diode
R42954 N42953 N42954 10
D42954 N42954 0 diode
R42955 N42954 N42955 10
D42955 N42955 0 diode
R42956 N42955 N42956 10
D42956 N42956 0 diode
R42957 N42956 N42957 10
D42957 N42957 0 diode
R42958 N42957 N42958 10
D42958 N42958 0 diode
R42959 N42958 N42959 10
D42959 N42959 0 diode
R42960 N42959 N42960 10
D42960 N42960 0 diode
R42961 N42960 N42961 10
D42961 N42961 0 diode
R42962 N42961 N42962 10
D42962 N42962 0 diode
R42963 N42962 N42963 10
D42963 N42963 0 diode
R42964 N42963 N42964 10
D42964 N42964 0 diode
R42965 N42964 N42965 10
D42965 N42965 0 diode
R42966 N42965 N42966 10
D42966 N42966 0 diode
R42967 N42966 N42967 10
D42967 N42967 0 diode
R42968 N42967 N42968 10
D42968 N42968 0 diode
R42969 N42968 N42969 10
D42969 N42969 0 diode
R42970 N42969 N42970 10
D42970 N42970 0 diode
R42971 N42970 N42971 10
D42971 N42971 0 diode
R42972 N42971 N42972 10
D42972 N42972 0 diode
R42973 N42972 N42973 10
D42973 N42973 0 diode
R42974 N42973 N42974 10
D42974 N42974 0 diode
R42975 N42974 N42975 10
D42975 N42975 0 diode
R42976 N42975 N42976 10
D42976 N42976 0 diode
R42977 N42976 N42977 10
D42977 N42977 0 diode
R42978 N42977 N42978 10
D42978 N42978 0 diode
R42979 N42978 N42979 10
D42979 N42979 0 diode
R42980 N42979 N42980 10
D42980 N42980 0 diode
R42981 N42980 N42981 10
D42981 N42981 0 diode
R42982 N42981 N42982 10
D42982 N42982 0 diode
R42983 N42982 N42983 10
D42983 N42983 0 diode
R42984 N42983 N42984 10
D42984 N42984 0 diode
R42985 N42984 N42985 10
D42985 N42985 0 diode
R42986 N42985 N42986 10
D42986 N42986 0 diode
R42987 N42986 N42987 10
D42987 N42987 0 diode
R42988 N42987 N42988 10
D42988 N42988 0 diode
R42989 N42988 N42989 10
D42989 N42989 0 diode
R42990 N42989 N42990 10
D42990 N42990 0 diode
R42991 N42990 N42991 10
D42991 N42991 0 diode
R42992 N42991 N42992 10
D42992 N42992 0 diode
R42993 N42992 N42993 10
D42993 N42993 0 diode
R42994 N42993 N42994 10
D42994 N42994 0 diode
R42995 N42994 N42995 10
D42995 N42995 0 diode
R42996 N42995 N42996 10
D42996 N42996 0 diode
R42997 N42996 N42997 10
D42997 N42997 0 diode
R42998 N42997 N42998 10
D42998 N42998 0 diode
R42999 N42998 N42999 10
D42999 N42999 0 diode
R43000 N42999 N43000 10
D43000 N43000 0 diode
R43001 N43000 N43001 10
D43001 N43001 0 diode
R43002 N43001 N43002 10
D43002 N43002 0 diode
R43003 N43002 N43003 10
D43003 N43003 0 diode
R43004 N43003 N43004 10
D43004 N43004 0 diode
R43005 N43004 N43005 10
D43005 N43005 0 diode
R43006 N43005 N43006 10
D43006 N43006 0 diode
R43007 N43006 N43007 10
D43007 N43007 0 diode
R43008 N43007 N43008 10
D43008 N43008 0 diode
R43009 N43008 N43009 10
D43009 N43009 0 diode
R43010 N43009 N43010 10
D43010 N43010 0 diode
R43011 N43010 N43011 10
D43011 N43011 0 diode
R43012 N43011 N43012 10
D43012 N43012 0 diode
R43013 N43012 N43013 10
D43013 N43013 0 diode
R43014 N43013 N43014 10
D43014 N43014 0 diode
R43015 N43014 N43015 10
D43015 N43015 0 diode
R43016 N43015 N43016 10
D43016 N43016 0 diode
R43017 N43016 N43017 10
D43017 N43017 0 diode
R43018 N43017 N43018 10
D43018 N43018 0 diode
R43019 N43018 N43019 10
D43019 N43019 0 diode
R43020 N43019 N43020 10
D43020 N43020 0 diode
R43021 N43020 N43021 10
D43021 N43021 0 diode
R43022 N43021 N43022 10
D43022 N43022 0 diode
R43023 N43022 N43023 10
D43023 N43023 0 diode
R43024 N43023 N43024 10
D43024 N43024 0 diode
R43025 N43024 N43025 10
D43025 N43025 0 diode
R43026 N43025 N43026 10
D43026 N43026 0 diode
R43027 N43026 N43027 10
D43027 N43027 0 diode
R43028 N43027 N43028 10
D43028 N43028 0 diode
R43029 N43028 N43029 10
D43029 N43029 0 diode
R43030 N43029 N43030 10
D43030 N43030 0 diode
R43031 N43030 N43031 10
D43031 N43031 0 diode
R43032 N43031 N43032 10
D43032 N43032 0 diode
R43033 N43032 N43033 10
D43033 N43033 0 diode
R43034 N43033 N43034 10
D43034 N43034 0 diode
R43035 N43034 N43035 10
D43035 N43035 0 diode
R43036 N43035 N43036 10
D43036 N43036 0 diode
R43037 N43036 N43037 10
D43037 N43037 0 diode
R43038 N43037 N43038 10
D43038 N43038 0 diode
R43039 N43038 N43039 10
D43039 N43039 0 diode
R43040 N43039 N43040 10
D43040 N43040 0 diode
R43041 N43040 N43041 10
D43041 N43041 0 diode
R43042 N43041 N43042 10
D43042 N43042 0 diode
R43043 N43042 N43043 10
D43043 N43043 0 diode
R43044 N43043 N43044 10
D43044 N43044 0 diode
R43045 N43044 N43045 10
D43045 N43045 0 diode
R43046 N43045 N43046 10
D43046 N43046 0 diode
R43047 N43046 N43047 10
D43047 N43047 0 diode
R43048 N43047 N43048 10
D43048 N43048 0 diode
R43049 N43048 N43049 10
D43049 N43049 0 diode
R43050 N43049 N43050 10
D43050 N43050 0 diode
R43051 N43050 N43051 10
D43051 N43051 0 diode
R43052 N43051 N43052 10
D43052 N43052 0 diode
R43053 N43052 N43053 10
D43053 N43053 0 diode
R43054 N43053 N43054 10
D43054 N43054 0 diode
R43055 N43054 N43055 10
D43055 N43055 0 diode
R43056 N43055 N43056 10
D43056 N43056 0 diode
R43057 N43056 N43057 10
D43057 N43057 0 diode
R43058 N43057 N43058 10
D43058 N43058 0 diode
R43059 N43058 N43059 10
D43059 N43059 0 diode
R43060 N43059 N43060 10
D43060 N43060 0 diode
R43061 N43060 N43061 10
D43061 N43061 0 diode
R43062 N43061 N43062 10
D43062 N43062 0 diode
R43063 N43062 N43063 10
D43063 N43063 0 diode
R43064 N43063 N43064 10
D43064 N43064 0 diode
R43065 N43064 N43065 10
D43065 N43065 0 diode
R43066 N43065 N43066 10
D43066 N43066 0 diode
R43067 N43066 N43067 10
D43067 N43067 0 diode
R43068 N43067 N43068 10
D43068 N43068 0 diode
R43069 N43068 N43069 10
D43069 N43069 0 diode
R43070 N43069 N43070 10
D43070 N43070 0 diode
R43071 N43070 N43071 10
D43071 N43071 0 diode
R43072 N43071 N43072 10
D43072 N43072 0 diode
R43073 N43072 N43073 10
D43073 N43073 0 diode
R43074 N43073 N43074 10
D43074 N43074 0 diode
R43075 N43074 N43075 10
D43075 N43075 0 diode
R43076 N43075 N43076 10
D43076 N43076 0 diode
R43077 N43076 N43077 10
D43077 N43077 0 diode
R43078 N43077 N43078 10
D43078 N43078 0 diode
R43079 N43078 N43079 10
D43079 N43079 0 diode
R43080 N43079 N43080 10
D43080 N43080 0 diode
R43081 N43080 N43081 10
D43081 N43081 0 diode
R43082 N43081 N43082 10
D43082 N43082 0 diode
R43083 N43082 N43083 10
D43083 N43083 0 diode
R43084 N43083 N43084 10
D43084 N43084 0 diode
R43085 N43084 N43085 10
D43085 N43085 0 diode
R43086 N43085 N43086 10
D43086 N43086 0 diode
R43087 N43086 N43087 10
D43087 N43087 0 diode
R43088 N43087 N43088 10
D43088 N43088 0 diode
R43089 N43088 N43089 10
D43089 N43089 0 diode
R43090 N43089 N43090 10
D43090 N43090 0 diode
R43091 N43090 N43091 10
D43091 N43091 0 diode
R43092 N43091 N43092 10
D43092 N43092 0 diode
R43093 N43092 N43093 10
D43093 N43093 0 diode
R43094 N43093 N43094 10
D43094 N43094 0 diode
R43095 N43094 N43095 10
D43095 N43095 0 diode
R43096 N43095 N43096 10
D43096 N43096 0 diode
R43097 N43096 N43097 10
D43097 N43097 0 diode
R43098 N43097 N43098 10
D43098 N43098 0 diode
R43099 N43098 N43099 10
D43099 N43099 0 diode
R43100 N43099 N43100 10
D43100 N43100 0 diode
R43101 N43100 N43101 10
D43101 N43101 0 diode
R43102 N43101 N43102 10
D43102 N43102 0 diode
R43103 N43102 N43103 10
D43103 N43103 0 diode
R43104 N43103 N43104 10
D43104 N43104 0 diode
R43105 N43104 N43105 10
D43105 N43105 0 diode
R43106 N43105 N43106 10
D43106 N43106 0 diode
R43107 N43106 N43107 10
D43107 N43107 0 diode
R43108 N43107 N43108 10
D43108 N43108 0 diode
R43109 N43108 N43109 10
D43109 N43109 0 diode
R43110 N43109 N43110 10
D43110 N43110 0 diode
R43111 N43110 N43111 10
D43111 N43111 0 diode
R43112 N43111 N43112 10
D43112 N43112 0 diode
R43113 N43112 N43113 10
D43113 N43113 0 diode
R43114 N43113 N43114 10
D43114 N43114 0 diode
R43115 N43114 N43115 10
D43115 N43115 0 diode
R43116 N43115 N43116 10
D43116 N43116 0 diode
R43117 N43116 N43117 10
D43117 N43117 0 diode
R43118 N43117 N43118 10
D43118 N43118 0 diode
R43119 N43118 N43119 10
D43119 N43119 0 diode
R43120 N43119 N43120 10
D43120 N43120 0 diode
R43121 N43120 N43121 10
D43121 N43121 0 diode
R43122 N43121 N43122 10
D43122 N43122 0 diode
R43123 N43122 N43123 10
D43123 N43123 0 diode
R43124 N43123 N43124 10
D43124 N43124 0 diode
R43125 N43124 N43125 10
D43125 N43125 0 diode
R43126 N43125 N43126 10
D43126 N43126 0 diode
R43127 N43126 N43127 10
D43127 N43127 0 diode
R43128 N43127 N43128 10
D43128 N43128 0 diode
R43129 N43128 N43129 10
D43129 N43129 0 diode
R43130 N43129 N43130 10
D43130 N43130 0 diode
R43131 N43130 N43131 10
D43131 N43131 0 diode
R43132 N43131 N43132 10
D43132 N43132 0 diode
R43133 N43132 N43133 10
D43133 N43133 0 diode
R43134 N43133 N43134 10
D43134 N43134 0 diode
R43135 N43134 N43135 10
D43135 N43135 0 diode
R43136 N43135 N43136 10
D43136 N43136 0 diode
R43137 N43136 N43137 10
D43137 N43137 0 diode
R43138 N43137 N43138 10
D43138 N43138 0 diode
R43139 N43138 N43139 10
D43139 N43139 0 diode
R43140 N43139 N43140 10
D43140 N43140 0 diode
R43141 N43140 N43141 10
D43141 N43141 0 diode
R43142 N43141 N43142 10
D43142 N43142 0 diode
R43143 N43142 N43143 10
D43143 N43143 0 diode
R43144 N43143 N43144 10
D43144 N43144 0 diode
R43145 N43144 N43145 10
D43145 N43145 0 diode
R43146 N43145 N43146 10
D43146 N43146 0 diode
R43147 N43146 N43147 10
D43147 N43147 0 diode
R43148 N43147 N43148 10
D43148 N43148 0 diode
R43149 N43148 N43149 10
D43149 N43149 0 diode
R43150 N43149 N43150 10
D43150 N43150 0 diode
R43151 N43150 N43151 10
D43151 N43151 0 diode
R43152 N43151 N43152 10
D43152 N43152 0 diode
R43153 N43152 N43153 10
D43153 N43153 0 diode
R43154 N43153 N43154 10
D43154 N43154 0 diode
R43155 N43154 N43155 10
D43155 N43155 0 diode
R43156 N43155 N43156 10
D43156 N43156 0 diode
R43157 N43156 N43157 10
D43157 N43157 0 diode
R43158 N43157 N43158 10
D43158 N43158 0 diode
R43159 N43158 N43159 10
D43159 N43159 0 diode
R43160 N43159 N43160 10
D43160 N43160 0 diode
R43161 N43160 N43161 10
D43161 N43161 0 diode
R43162 N43161 N43162 10
D43162 N43162 0 diode
R43163 N43162 N43163 10
D43163 N43163 0 diode
R43164 N43163 N43164 10
D43164 N43164 0 diode
R43165 N43164 N43165 10
D43165 N43165 0 diode
R43166 N43165 N43166 10
D43166 N43166 0 diode
R43167 N43166 N43167 10
D43167 N43167 0 diode
R43168 N43167 N43168 10
D43168 N43168 0 diode
R43169 N43168 N43169 10
D43169 N43169 0 diode
R43170 N43169 N43170 10
D43170 N43170 0 diode
R43171 N43170 N43171 10
D43171 N43171 0 diode
R43172 N43171 N43172 10
D43172 N43172 0 diode
R43173 N43172 N43173 10
D43173 N43173 0 diode
R43174 N43173 N43174 10
D43174 N43174 0 diode
R43175 N43174 N43175 10
D43175 N43175 0 diode
R43176 N43175 N43176 10
D43176 N43176 0 diode
R43177 N43176 N43177 10
D43177 N43177 0 diode
R43178 N43177 N43178 10
D43178 N43178 0 diode
R43179 N43178 N43179 10
D43179 N43179 0 diode
R43180 N43179 N43180 10
D43180 N43180 0 diode
R43181 N43180 N43181 10
D43181 N43181 0 diode
R43182 N43181 N43182 10
D43182 N43182 0 diode
R43183 N43182 N43183 10
D43183 N43183 0 diode
R43184 N43183 N43184 10
D43184 N43184 0 diode
R43185 N43184 N43185 10
D43185 N43185 0 diode
R43186 N43185 N43186 10
D43186 N43186 0 diode
R43187 N43186 N43187 10
D43187 N43187 0 diode
R43188 N43187 N43188 10
D43188 N43188 0 diode
R43189 N43188 N43189 10
D43189 N43189 0 diode
R43190 N43189 N43190 10
D43190 N43190 0 diode
R43191 N43190 N43191 10
D43191 N43191 0 diode
R43192 N43191 N43192 10
D43192 N43192 0 diode
R43193 N43192 N43193 10
D43193 N43193 0 diode
R43194 N43193 N43194 10
D43194 N43194 0 diode
R43195 N43194 N43195 10
D43195 N43195 0 diode
R43196 N43195 N43196 10
D43196 N43196 0 diode
R43197 N43196 N43197 10
D43197 N43197 0 diode
R43198 N43197 N43198 10
D43198 N43198 0 diode
R43199 N43198 N43199 10
D43199 N43199 0 diode
R43200 N43199 N43200 10
D43200 N43200 0 diode
R43201 N43200 N43201 10
D43201 N43201 0 diode
R43202 N43201 N43202 10
D43202 N43202 0 diode
R43203 N43202 N43203 10
D43203 N43203 0 diode
R43204 N43203 N43204 10
D43204 N43204 0 diode
R43205 N43204 N43205 10
D43205 N43205 0 diode
R43206 N43205 N43206 10
D43206 N43206 0 diode
R43207 N43206 N43207 10
D43207 N43207 0 diode
R43208 N43207 N43208 10
D43208 N43208 0 diode
R43209 N43208 N43209 10
D43209 N43209 0 diode
R43210 N43209 N43210 10
D43210 N43210 0 diode
R43211 N43210 N43211 10
D43211 N43211 0 diode
R43212 N43211 N43212 10
D43212 N43212 0 diode
R43213 N43212 N43213 10
D43213 N43213 0 diode
R43214 N43213 N43214 10
D43214 N43214 0 diode
R43215 N43214 N43215 10
D43215 N43215 0 diode
R43216 N43215 N43216 10
D43216 N43216 0 diode
R43217 N43216 N43217 10
D43217 N43217 0 diode
R43218 N43217 N43218 10
D43218 N43218 0 diode
R43219 N43218 N43219 10
D43219 N43219 0 diode
R43220 N43219 N43220 10
D43220 N43220 0 diode
R43221 N43220 N43221 10
D43221 N43221 0 diode
R43222 N43221 N43222 10
D43222 N43222 0 diode
R43223 N43222 N43223 10
D43223 N43223 0 diode
R43224 N43223 N43224 10
D43224 N43224 0 diode
R43225 N43224 N43225 10
D43225 N43225 0 diode
R43226 N43225 N43226 10
D43226 N43226 0 diode
R43227 N43226 N43227 10
D43227 N43227 0 diode
R43228 N43227 N43228 10
D43228 N43228 0 diode
R43229 N43228 N43229 10
D43229 N43229 0 diode
R43230 N43229 N43230 10
D43230 N43230 0 diode
R43231 N43230 N43231 10
D43231 N43231 0 diode
R43232 N43231 N43232 10
D43232 N43232 0 diode
R43233 N43232 N43233 10
D43233 N43233 0 diode
R43234 N43233 N43234 10
D43234 N43234 0 diode
R43235 N43234 N43235 10
D43235 N43235 0 diode
R43236 N43235 N43236 10
D43236 N43236 0 diode
R43237 N43236 N43237 10
D43237 N43237 0 diode
R43238 N43237 N43238 10
D43238 N43238 0 diode
R43239 N43238 N43239 10
D43239 N43239 0 diode
R43240 N43239 N43240 10
D43240 N43240 0 diode
R43241 N43240 N43241 10
D43241 N43241 0 diode
R43242 N43241 N43242 10
D43242 N43242 0 diode
R43243 N43242 N43243 10
D43243 N43243 0 diode
R43244 N43243 N43244 10
D43244 N43244 0 diode
R43245 N43244 N43245 10
D43245 N43245 0 diode
R43246 N43245 N43246 10
D43246 N43246 0 diode
R43247 N43246 N43247 10
D43247 N43247 0 diode
R43248 N43247 N43248 10
D43248 N43248 0 diode
R43249 N43248 N43249 10
D43249 N43249 0 diode
R43250 N43249 N43250 10
D43250 N43250 0 diode
R43251 N43250 N43251 10
D43251 N43251 0 diode
R43252 N43251 N43252 10
D43252 N43252 0 diode
R43253 N43252 N43253 10
D43253 N43253 0 diode
R43254 N43253 N43254 10
D43254 N43254 0 diode
R43255 N43254 N43255 10
D43255 N43255 0 diode
R43256 N43255 N43256 10
D43256 N43256 0 diode
R43257 N43256 N43257 10
D43257 N43257 0 diode
R43258 N43257 N43258 10
D43258 N43258 0 diode
R43259 N43258 N43259 10
D43259 N43259 0 diode
R43260 N43259 N43260 10
D43260 N43260 0 diode
R43261 N43260 N43261 10
D43261 N43261 0 diode
R43262 N43261 N43262 10
D43262 N43262 0 diode
R43263 N43262 N43263 10
D43263 N43263 0 diode
R43264 N43263 N43264 10
D43264 N43264 0 diode
R43265 N43264 N43265 10
D43265 N43265 0 diode
R43266 N43265 N43266 10
D43266 N43266 0 diode
R43267 N43266 N43267 10
D43267 N43267 0 diode
R43268 N43267 N43268 10
D43268 N43268 0 diode
R43269 N43268 N43269 10
D43269 N43269 0 diode
R43270 N43269 N43270 10
D43270 N43270 0 diode
R43271 N43270 N43271 10
D43271 N43271 0 diode
R43272 N43271 N43272 10
D43272 N43272 0 diode
R43273 N43272 N43273 10
D43273 N43273 0 diode
R43274 N43273 N43274 10
D43274 N43274 0 diode
R43275 N43274 N43275 10
D43275 N43275 0 diode
R43276 N43275 N43276 10
D43276 N43276 0 diode
R43277 N43276 N43277 10
D43277 N43277 0 diode
R43278 N43277 N43278 10
D43278 N43278 0 diode
R43279 N43278 N43279 10
D43279 N43279 0 diode
R43280 N43279 N43280 10
D43280 N43280 0 diode
R43281 N43280 N43281 10
D43281 N43281 0 diode
R43282 N43281 N43282 10
D43282 N43282 0 diode
R43283 N43282 N43283 10
D43283 N43283 0 diode
R43284 N43283 N43284 10
D43284 N43284 0 diode
R43285 N43284 N43285 10
D43285 N43285 0 diode
R43286 N43285 N43286 10
D43286 N43286 0 diode
R43287 N43286 N43287 10
D43287 N43287 0 diode
R43288 N43287 N43288 10
D43288 N43288 0 diode
R43289 N43288 N43289 10
D43289 N43289 0 diode
R43290 N43289 N43290 10
D43290 N43290 0 diode
R43291 N43290 N43291 10
D43291 N43291 0 diode
R43292 N43291 N43292 10
D43292 N43292 0 diode
R43293 N43292 N43293 10
D43293 N43293 0 diode
R43294 N43293 N43294 10
D43294 N43294 0 diode
R43295 N43294 N43295 10
D43295 N43295 0 diode
R43296 N43295 N43296 10
D43296 N43296 0 diode
R43297 N43296 N43297 10
D43297 N43297 0 diode
R43298 N43297 N43298 10
D43298 N43298 0 diode
R43299 N43298 N43299 10
D43299 N43299 0 diode
R43300 N43299 N43300 10
D43300 N43300 0 diode
R43301 N43300 N43301 10
D43301 N43301 0 diode
R43302 N43301 N43302 10
D43302 N43302 0 diode
R43303 N43302 N43303 10
D43303 N43303 0 diode
R43304 N43303 N43304 10
D43304 N43304 0 diode
R43305 N43304 N43305 10
D43305 N43305 0 diode
R43306 N43305 N43306 10
D43306 N43306 0 diode
R43307 N43306 N43307 10
D43307 N43307 0 diode
R43308 N43307 N43308 10
D43308 N43308 0 diode
R43309 N43308 N43309 10
D43309 N43309 0 diode
R43310 N43309 N43310 10
D43310 N43310 0 diode
R43311 N43310 N43311 10
D43311 N43311 0 diode
R43312 N43311 N43312 10
D43312 N43312 0 diode
R43313 N43312 N43313 10
D43313 N43313 0 diode
R43314 N43313 N43314 10
D43314 N43314 0 diode
R43315 N43314 N43315 10
D43315 N43315 0 diode
R43316 N43315 N43316 10
D43316 N43316 0 diode
R43317 N43316 N43317 10
D43317 N43317 0 diode
R43318 N43317 N43318 10
D43318 N43318 0 diode
R43319 N43318 N43319 10
D43319 N43319 0 diode
R43320 N43319 N43320 10
D43320 N43320 0 diode
R43321 N43320 N43321 10
D43321 N43321 0 diode
R43322 N43321 N43322 10
D43322 N43322 0 diode
R43323 N43322 N43323 10
D43323 N43323 0 diode
R43324 N43323 N43324 10
D43324 N43324 0 diode
R43325 N43324 N43325 10
D43325 N43325 0 diode
R43326 N43325 N43326 10
D43326 N43326 0 diode
R43327 N43326 N43327 10
D43327 N43327 0 diode
R43328 N43327 N43328 10
D43328 N43328 0 diode
R43329 N43328 N43329 10
D43329 N43329 0 diode
R43330 N43329 N43330 10
D43330 N43330 0 diode
R43331 N43330 N43331 10
D43331 N43331 0 diode
R43332 N43331 N43332 10
D43332 N43332 0 diode
R43333 N43332 N43333 10
D43333 N43333 0 diode
R43334 N43333 N43334 10
D43334 N43334 0 diode
R43335 N43334 N43335 10
D43335 N43335 0 diode
R43336 N43335 N43336 10
D43336 N43336 0 diode
R43337 N43336 N43337 10
D43337 N43337 0 diode
R43338 N43337 N43338 10
D43338 N43338 0 diode
R43339 N43338 N43339 10
D43339 N43339 0 diode
R43340 N43339 N43340 10
D43340 N43340 0 diode
R43341 N43340 N43341 10
D43341 N43341 0 diode
R43342 N43341 N43342 10
D43342 N43342 0 diode
R43343 N43342 N43343 10
D43343 N43343 0 diode
R43344 N43343 N43344 10
D43344 N43344 0 diode
R43345 N43344 N43345 10
D43345 N43345 0 diode
R43346 N43345 N43346 10
D43346 N43346 0 diode
R43347 N43346 N43347 10
D43347 N43347 0 diode
R43348 N43347 N43348 10
D43348 N43348 0 diode
R43349 N43348 N43349 10
D43349 N43349 0 diode
R43350 N43349 N43350 10
D43350 N43350 0 diode
R43351 N43350 N43351 10
D43351 N43351 0 diode
R43352 N43351 N43352 10
D43352 N43352 0 diode
R43353 N43352 N43353 10
D43353 N43353 0 diode
R43354 N43353 N43354 10
D43354 N43354 0 diode
R43355 N43354 N43355 10
D43355 N43355 0 diode
R43356 N43355 N43356 10
D43356 N43356 0 diode
R43357 N43356 N43357 10
D43357 N43357 0 diode
R43358 N43357 N43358 10
D43358 N43358 0 diode
R43359 N43358 N43359 10
D43359 N43359 0 diode
R43360 N43359 N43360 10
D43360 N43360 0 diode
R43361 N43360 N43361 10
D43361 N43361 0 diode
R43362 N43361 N43362 10
D43362 N43362 0 diode
R43363 N43362 N43363 10
D43363 N43363 0 diode
R43364 N43363 N43364 10
D43364 N43364 0 diode
R43365 N43364 N43365 10
D43365 N43365 0 diode
R43366 N43365 N43366 10
D43366 N43366 0 diode
R43367 N43366 N43367 10
D43367 N43367 0 diode
R43368 N43367 N43368 10
D43368 N43368 0 diode
R43369 N43368 N43369 10
D43369 N43369 0 diode
R43370 N43369 N43370 10
D43370 N43370 0 diode
R43371 N43370 N43371 10
D43371 N43371 0 diode
R43372 N43371 N43372 10
D43372 N43372 0 diode
R43373 N43372 N43373 10
D43373 N43373 0 diode
R43374 N43373 N43374 10
D43374 N43374 0 diode
R43375 N43374 N43375 10
D43375 N43375 0 diode
R43376 N43375 N43376 10
D43376 N43376 0 diode
R43377 N43376 N43377 10
D43377 N43377 0 diode
R43378 N43377 N43378 10
D43378 N43378 0 diode
R43379 N43378 N43379 10
D43379 N43379 0 diode
R43380 N43379 N43380 10
D43380 N43380 0 diode
R43381 N43380 N43381 10
D43381 N43381 0 diode
R43382 N43381 N43382 10
D43382 N43382 0 diode
R43383 N43382 N43383 10
D43383 N43383 0 diode
R43384 N43383 N43384 10
D43384 N43384 0 diode
R43385 N43384 N43385 10
D43385 N43385 0 diode
R43386 N43385 N43386 10
D43386 N43386 0 diode
R43387 N43386 N43387 10
D43387 N43387 0 diode
R43388 N43387 N43388 10
D43388 N43388 0 diode
R43389 N43388 N43389 10
D43389 N43389 0 diode
R43390 N43389 N43390 10
D43390 N43390 0 diode
R43391 N43390 N43391 10
D43391 N43391 0 diode
R43392 N43391 N43392 10
D43392 N43392 0 diode
R43393 N43392 N43393 10
D43393 N43393 0 diode
R43394 N43393 N43394 10
D43394 N43394 0 diode
R43395 N43394 N43395 10
D43395 N43395 0 diode
R43396 N43395 N43396 10
D43396 N43396 0 diode
R43397 N43396 N43397 10
D43397 N43397 0 diode
R43398 N43397 N43398 10
D43398 N43398 0 diode
R43399 N43398 N43399 10
D43399 N43399 0 diode
R43400 N43399 N43400 10
D43400 N43400 0 diode
R43401 N43400 N43401 10
D43401 N43401 0 diode
R43402 N43401 N43402 10
D43402 N43402 0 diode
R43403 N43402 N43403 10
D43403 N43403 0 diode
R43404 N43403 N43404 10
D43404 N43404 0 diode
R43405 N43404 N43405 10
D43405 N43405 0 diode
R43406 N43405 N43406 10
D43406 N43406 0 diode
R43407 N43406 N43407 10
D43407 N43407 0 diode
R43408 N43407 N43408 10
D43408 N43408 0 diode
R43409 N43408 N43409 10
D43409 N43409 0 diode
R43410 N43409 N43410 10
D43410 N43410 0 diode
R43411 N43410 N43411 10
D43411 N43411 0 diode
R43412 N43411 N43412 10
D43412 N43412 0 diode
R43413 N43412 N43413 10
D43413 N43413 0 diode
R43414 N43413 N43414 10
D43414 N43414 0 diode
R43415 N43414 N43415 10
D43415 N43415 0 diode
R43416 N43415 N43416 10
D43416 N43416 0 diode
R43417 N43416 N43417 10
D43417 N43417 0 diode
R43418 N43417 N43418 10
D43418 N43418 0 diode
R43419 N43418 N43419 10
D43419 N43419 0 diode
R43420 N43419 N43420 10
D43420 N43420 0 diode
R43421 N43420 N43421 10
D43421 N43421 0 diode
R43422 N43421 N43422 10
D43422 N43422 0 diode
R43423 N43422 N43423 10
D43423 N43423 0 diode
R43424 N43423 N43424 10
D43424 N43424 0 diode
R43425 N43424 N43425 10
D43425 N43425 0 diode
R43426 N43425 N43426 10
D43426 N43426 0 diode
R43427 N43426 N43427 10
D43427 N43427 0 diode
R43428 N43427 N43428 10
D43428 N43428 0 diode
R43429 N43428 N43429 10
D43429 N43429 0 diode
R43430 N43429 N43430 10
D43430 N43430 0 diode
R43431 N43430 N43431 10
D43431 N43431 0 diode
R43432 N43431 N43432 10
D43432 N43432 0 diode
R43433 N43432 N43433 10
D43433 N43433 0 diode
R43434 N43433 N43434 10
D43434 N43434 0 diode
R43435 N43434 N43435 10
D43435 N43435 0 diode
R43436 N43435 N43436 10
D43436 N43436 0 diode
R43437 N43436 N43437 10
D43437 N43437 0 diode
R43438 N43437 N43438 10
D43438 N43438 0 diode
R43439 N43438 N43439 10
D43439 N43439 0 diode
R43440 N43439 N43440 10
D43440 N43440 0 diode
R43441 N43440 N43441 10
D43441 N43441 0 diode
R43442 N43441 N43442 10
D43442 N43442 0 diode
R43443 N43442 N43443 10
D43443 N43443 0 diode
R43444 N43443 N43444 10
D43444 N43444 0 diode
R43445 N43444 N43445 10
D43445 N43445 0 diode
R43446 N43445 N43446 10
D43446 N43446 0 diode
R43447 N43446 N43447 10
D43447 N43447 0 diode
R43448 N43447 N43448 10
D43448 N43448 0 diode
R43449 N43448 N43449 10
D43449 N43449 0 diode
R43450 N43449 N43450 10
D43450 N43450 0 diode
R43451 N43450 N43451 10
D43451 N43451 0 diode
R43452 N43451 N43452 10
D43452 N43452 0 diode
R43453 N43452 N43453 10
D43453 N43453 0 diode
R43454 N43453 N43454 10
D43454 N43454 0 diode
R43455 N43454 N43455 10
D43455 N43455 0 diode
R43456 N43455 N43456 10
D43456 N43456 0 diode
R43457 N43456 N43457 10
D43457 N43457 0 diode
R43458 N43457 N43458 10
D43458 N43458 0 diode
R43459 N43458 N43459 10
D43459 N43459 0 diode
R43460 N43459 N43460 10
D43460 N43460 0 diode
R43461 N43460 N43461 10
D43461 N43461 0 diode
R43462 N43461 N43462 10
D43462 N43462 0 diode
R43463 N43462 N43463 10
D43463 N43463 0 diode
R43464 N43463 N43464 10
D43464 N43464 0 diode
R43465 N43464 N43465 10
D43465 N43465 0 diode
R43466 N43465 N43466 10
D43466 N43466 0 diode
R43467 N43466 N43467 10
D43467 N43467 0 diode
R43468 N43467 N43468 10
D43468 N43468 0 diode
R43469 N43468 N43469 10
D43469 N43469 0 diode
R43470 N43469 N43470 10
D43470 N43470 0 diode
R43471 N43470 N43471 10
D43471 N43471 0 diode
R43472 N43471 N43472 10
D43472 N43472 0 diode
R43473 N43472 N43473 10
D43473 N43473 0 diode
R43474 N43473 N43474 10
D43474 N43474 0 diode
R43475 N43474 N43475 10
D43475 N43475 0 diode
R43476 N43475 N43476 10
D43476 N43476 0 diode
R43477 N43476 N43477 10
D43477 N43477 0 diode
R43478 N43477 N43478 10
D43478 N43478 0 diode
R43479 N43478 N43479 10
D43479 N43479 0 diode
R43480 N43479 N43480 10
D43480 N43480 0 diode
R43481 N43480 N43481 10
D43481 N43481 0 diode
R43482 N43481 N43482 10
D43482 N43482 0 diode
R43483 N43482 N43483 10
D43483 N43483 0 diode
R43484 N43483 N43484 10
D43484 N43484 0 diode
R43485 N43484 N43485 10
D43485 N43485 0 diode
R43486 N43485 N43486 10
D43486 N43486 0 diode
R43487 N43486 N43487 10
D43487 N43487 0 diode
R43488 N43487 N43488 10
D43488 N43488 0 diode
R43489 N43488 N43489 10
D43489 N43489 0 diode
R43490 N43489 N43490 10
D43490 N43490 0 diode
R43491 N43490 N43491 10
D43491 N43491 0 diode
R43492 N43491 N43492 10
D43492 N43492 0 diode
R43493 N43492 N43493 10
D43493 N43493 0 diode
R43494 N43493 N43494 10
D43494 N43494 0 diode
R43495 N43494 N43495 10
D43495 N43495 0 diode
R43496 N43495 N43496 10
D43496 N43496 0 diode
R43497 N43496 N43497 10
D43497 N43497 0 diode
R43498 N43497 N43498 10
D43498 N43498 0 diode
R43499 N43498 N43499 10
D43499 N43499 0 diode
R43500 N43499 N43500 10
D43500 N43500 0 diode
R43501 N43500 N43501 10
D43501 N43501 0 diode
R43502 N43501 N43502 10
D43502 N43502 0 diode
R43503 N43502 N43503 10
D43503 N43503 0 diode
R43504 N43503 N43504 10
D43504 N43504 0 diode
R43505 N43504 N43505 10
D43505 N43505 0 diode
R43506 N43505 N43506 10
D43506 N43506 0 diode
R43507 N43506 N43507 10
D43507 N43507 0 diode
R43508 N43507 N43508 10
D43508 N43508 0 diode
R43509 N43508 N43509 10
D43509 N43509 0 diode
R43510 N43509 N43510 10
D43510 N43510 0 diode
R43511 N43510 N43511 10
D43511 N43511 0 diode
R43512 N43511 N43512 10
D43512 N43512 0 diode
R43513 N43512 N43513 10
D43513 N43513 0 diode
R43514 N43513 N43514 10
D43514 N43514 0 diode
R43515 N43514 N43515 10
D43515 N43515 0 diode
R43516 N43515 N43516 10
D43516 N43516 0 diode
R43517 N43516 N43517 10
D43517 N43517 0 diode
R43518 N43517 N43518 10
D43518 N43518 0 diode
R43519 N43518 N43519 10
D43519 N43519 0 diode
R43520 N43519 N43520 10
D43520 N43520 0 diode
R43521 N43520 N43521 10
D43521 N43521 0 diode
R43522 N43521 N43522 10
D43522 N43522 0 diode
R43523 N43522 N43523 10
D43523 N43523 0 diode
R43524 N43523 N43524 10
D43524 N43524 0 diode
R43525 N43524 N43525 10
D43525 N43525 0 diode
R43526 N43525 N43526 10
D43526 N43526 0 diode
R43527 N43526 N43527 10
D43527 N43527 0 diode
R43528 N43527 N43528 10
D43528 N43528 0 diode
R43529 N43528 N43529 10
D43529 N43529 0 diode
R43530 N43529 N43530 10
D43530 N43530 0 diode
R43531 N43530 N43531 10
D43531 N43531 0 diode
R43532 N43531 N43532 10
D43532 N43532 0 diode
R43533 N43532 N43533 10
D43533 N43533 0 diode
R43534 N43533 N43534 10
D43534 N43534 0 diode
R43535 N43534 N43535 10
D43535 N43535 0 diode
R43536 N43535 N43536 10
D43536 N43536 0 diode
R43537 N43536 N43537 10
D43537 N43537 0 diode
R43538 N43537 N43538 10
D43538 N43538 0 diode
R43539 N43538 N43539 10
D43539 N43539 0 diode
R43540 N43539 N43540 10
D43540 N43540 0 diode
R43541 N43540 N43541 10
D43541 N43541 0 diode
R43542 N43541 N43542 10
D43542 N43542 0 diode
R43543 N43542 N43543 10
D43543 N43543 0 diode
R43544 N43543 N43544 10
D43544 N43544 0 diode
R43545 N43544 N43545 10
D43545 N43545 0 diode
R43546 N43545 N43546 10
D43546 N43546 0 diode
R43547 N43546 N43547 10
D43547 N43547 0 diode
R43548 N43547 N43548 10
D43548 N43548 0 diode
R43549 N43548 N43549 10
D43549 N43549 0 diode
R43550 N43549 N43550 10
D43550 N43550 0 diode
R43551 N43550 N43551 10
D43551 N43551 0 diode
R43552 N43551 N43552 10
D43552 N43552 0 diode
R43553 N43552 N43553 10
D43553 N43553 0 diode
R43554 N43553 N43554 10
D43554 N43554 0 diode
R43555 N43554 N43555 10
D43555 N43555 0 diode
R43556 N43555 N43556 10
D43556 N43556 0 diode
R43557 N43556 N43557 10
D43557 N43557 0 diode
R43558 N43557 N43558 10
D43558 N43558 0 diode
R43559 N43558 N43559 10
D43559 N43559 0 diode
R43560 N43559 N43560 10
D43560 N43560 0 diode
R43561 N43560 N43561 10
D43561 N43561 0 diode
R43562 N43561 N43562 10
D43562 N43562 0 diode
R43563 N43562 N43563 10
D43563 N43563 0 diode
R43564 N43563 N43564 10
D43564 N43564 0 diode
R43565 N43564 N43565 10
D43565 N43565 0 diode
R43566 N43565 N43566 10
D43566 N43566 0 diode
R43567 N43566 N43567 10
D43567 N43567 0 diode
R43568 N43567 N43568 10
D43568 N43568 0 diode
R43569 N43568 N43569 10
D43569 N43569 0 diode
R43570 N43569 N43570 10
D43570 N43570 0 diode
R43571 N43570 N43571 10
D43571 N43571 0 diode
R43572 N43571 N43572 10
D43572 N43572 0 diode
R43573 N43572 N43573 10
D43573 N43573 0 diode
R43574 N43573 N43574 10
D43574 N43574 0 diode
R43575 N43574 N43575 10
D43575 N43575 0 diode
R43576 N43575 N43576 10
D43576 N43576 0 diode
R43577 N43576 N43577 10
D43577 N43577 0 diode
R43578 N43577 N43578 10
D43578 N43578 0 diode
R43579 N43578 N43579 10
D43579 N43579 0 diode
R43580 N43579 N43580 10
D43580 N43580 0 diode
R43581 N43580 N43581 10
D43581 N43581 0 diode
R43582 N43581 N43582 10
D43582 N43582 0 diode
R43583 N43582 N43583 10
D43583 N43583 0 diode
R43584 N43583 N43584 10
D43584 N43584 0 diode
R43585 N43584 N43585 10
D43585 N43585 0 diode
R43586 N43585 N43586 10
D43586 N43586 0 diode
R43587 N43586 N43587 10
D43587 N43587 0 diode
R43588 N43587 N43588 10
D43588 N43588 0 diode
R43589 N43588 N43589 10
D43589 N43589 0 diode
R43590 N43589 N43590 10
D43590 N43590 0 diode
R43591 N43590 N43591 10
D43591 N43591 0 diode
R43592 N43591 N43592 10
D43592 N43592 0 diode
R43593 N43592 N43593 10
D43593 N43593 0 diode
R43594 N43593 N43594 10
D43594 N43594 0 diode
R43595 N43594 N43595 10
D43595 N43595 0 diode
R43596 N43595 N43596 10
D43596 N43596 0 diode
R43597 N43596 N43597 10
D43597 N43597 0 diode
R43598 N43597 N43598 10
D43598 N43598 0 diode
R43599 N43598 N43599 10
D43599 N43599 0 diode
R43600 N43599 N43600 10
D43600 N43600 0 diode
R43601 N43600 N43601 10
D43601 N43601 0 diode
R43602 N43601 N43602 10
D43602 N43602 0 diode
R43603 N43602 N43603 10
D43603 N43603 0 diode
R43604 N43603 N43604 10
D43604 N43604 0 diode
R43605 N43604 N43605 10
D43605 N43605 0 diode
R43606 N43605 N43606 10
D43606 N43606 0 diode
R43607 N43606 N43607 10
D43607 N43607 0 diode
R43608 N43607 N43608 10
D43608 N43608 0 diode
R43609 N43608 N43609 10
D43609 N43609 0 diode
R43610 N43609 N43610 10
D43610 N43610 0 diode
R43611 N43610 N43611 10
D43611 N43611 0 diode
R43612 N43611 N43612 10
D43612 N43612 0 diode
R43613 N43612 N43613 10
D43613 N43613 0 diode
R43614 N43613 N43614 10
D43614 N43614 0 diode
R43615 N43614 N43615 10
D43615 N43615 0 diode
R43616 N43615 N43616 10
D43616 N43616 0 diode
R43617 N43616 N43617 10
D43617 N43617 0 diode
R43618 N43617 N43618 10
D43618 N43618 0 diode
R43619 N43618 N43619 10
D43619 N43619 0 diode
R43620 N43619 N43620 10
D43620 N43620 0 diode
R43621 N43620 N43621 10
D43621 N43621 0 diode
R43622 N43621 N43622 10
D43622 N43622 0 diode
R43623 N43622 N43623 10
D43623 N43623 0 diode
R43624 N43623 N43624 10
D43624 N43624 0 diode
R43625 N43624 N43625 10
D43625 N43625 0 diode
R43626 N43625 N43626 10
D43626 N43626 0 diode
R43627 N43626 N43627 10
D43627 N43627 0 diode
R43628 N43627 N43628 10
D43628 N43628 0 diode
R43629 N43628 N43629 10
D43629 N43629 0 diode
R43630 N43629 N43630 10
D43630 N43630 0 diode
R43631 N43630 N43631 10
D43631 N43631 0 diode
R43632 N43631 N43632 10
D43632 N43632 0 diode
R43633 N43632 N43633 10
D43633 N43633 0 diode
R43634 N43633 N43634 10
D43634 N43634 0 diode
R43635 N43634 N43635 10
D43635 N43635 0 diode
R43636 N43635 N43636 10
D43636 N43636 0 diode
R43637 N43636 N43637 10
D43637 N43637 0 diode
R43638 N43637 N43638 10
D43638 N43638 0 diode
R43639 N43638 N43639 10
D43639 N43639 0 diode
R43640 N43639 N43640 10
D43640 N43640 0 diode
R43641 N43640 N43641 10
D43641 N43641 0 diode
R43642 N43641 N43642 10
D43642 N43642 0 diode
R43643 N43642 N43643 10
D43643 N43643 0 diode
R43644 N43643 N43644 10
D43644 N43644 0 diode
R43645 N43644 N43645 10
D43645 N43645 0 diode
R43646 N43645 N43646 10
D43646 N43646 0 diode
R43647 N43646 N43647 10
D43647 N43647 0 diode
R43648 N43647 N43648 10
D43648 N43648 0 diode
R43649 N43648 N43649 10
D43649 N43649 0 diode
R43650 N43649 N43650 10
D43650 N43650 0 diode
R43651 N43650 N43651 10
D43651 N43651 0 diode
R43652 N43651 N43652 10
D43652 N43652 0 diode
R43653 N43652 N43653 10
D43653 N43653 0 diode
R43654 N43653 N43654 10
D43654 N43654 0 diode
R43655 N43654 N43655 10
D43655 N43655 0 diode
R43656 N43655 N43656 10
D43656 N43656 0 diode
R43657 N43656 N43657 10
D43657 N43657 0 diode
R43658 N43657 N43658 10
D43658 N43658 0 diode
R43659 N43658 N43659 10
D43659 N43659 0 diode
R43660 N43659 N43660 10
D43660 N43660 0 diode
R43661 N43660 N43661 10
D43661 N43661 0 diode
R43662 N43661 N43662 10
D43662 N43662 0 diode
R43663 N43662 N43663 10
D43663 N43663 0 diode
R43664 N43663 N43664 10
D43664 N43664 0 diode
R43665 N43664 N43665 10
D43665 N43665 0 diode
R43666 N43665 N43666 10
D43666 N43666 0 diode
R43667 N43666 N43667 10
D43667 N43667 0 diode
R43668 N43667 N43668 10
D43668 N43668 0 diode
R43669 N43668 N43669 10
D43669 N43669 0 diode
R43670 N43669 N43670 10
D43670 N43670 0 diode
R43671 N43670 N43671 10
D43671 N43671 0 diode
R43672 N43671 N43672 10
D43672 N43672 0 diode
R43673 N43672 N43673 10
D43673 N43673 0 diode
R43674 N43673 N43674 10
D43674 N43674 0 diode
R43675 N43674 N43675 10
D43675 N43675 0 diode
R43676 N43675 N43676 10
D43676 N43676 0 diode
R43677 N43676 N43677 10
D43677 N43677 0 diode
R43678 N43677 N43678 10
D43678 N43678 0 diode
R43679 N43678 N43679 10
D43679 N43679 0 diode
R43680 N43679 N43680 10
D43680 N43680 0 diode
R43681 N43680 N43681 10
D43681 N43681 0 diode
R43682 N43681 N43682 10
D43682 N43682 0 diode
R43683 N43682 N43683 10
D43683 N43683 0 diode
R43684 N43683 N43684 10
D43684 N43684 0 diode
R43685 N43684 N43685 10
D43685 N43685 0 diode
R43686 N43685 N43686 10
D43686 N43686 0 diode
R43687 N43686 N43687 10
D43687 N43687 0 diode
R43688 N43687 N43688 10
D43688 N43688 0 diode
R43689 N43688 N43689 10
D43689 N43689 0 diode
R43690 N43689 N43690 10
D43690 N43690 0 diode
R43691 N43690 N43691 10
D43691 N43691 0 diode
R43692 N43691 N43692 10
D43692 N43692 0 diode
R43693 N43692 N43693 10
D43693 N43693 0 diode
R43694 N43693 N43694 10
D43694 N43694 0 diode
R43695 N43694 N43695 10
D43695 N43695 0 diode
R43696 N43695 N43696 10
D43696 N43696 0 diode
R43697 N43696 N43697 10
D43697 N43697 0 diode
R43698 N43697 N43698 10
D43698 N43698 0 diode
R43699 N43698 N43699 10
D43699 N43699 0 diode
R43700 N43699 N43700 10
D43700 N43700 0 diode
R43701 N43700 N43701 10
D43701 N43701 0 diode
R43702 N43701 N43702 10
D43702 N43702 0 diode
R43703 N43702 N43703 10
D43703 N43703 0 diode
R43704 N43703 N43704 10
D43704 N43704 0 diode
R43705 N43704 N43705 10
D43705 N43705 0 diode
R43706 N43705 N43706 10
D43706 N43706 0 diode
R43707 N43706 N43707 10
D43707 N43707 0 diode
R43708 N43707 N43708 10
D43708 N43708 0 diode
R43709 N43708 N43709 10
D43709 N43709 0 diode
R43710 N43709 N43710 10
D43710 N43710 0 diode
R43711 N43710 N43711 10
D43711 N43711 0 diode
R43712 N43711 N43712 10
D43712 N43712 0 diode
R43713 N43712 N43713 10
D43713 N43713 0 diode
R43714 N43713 N43714 10
D43714 N43714 0 diode
R43715 N43714 N43715 10
D43715 N43715 0 diode
R43716 N43715 N43716 10
D43716 N43716 0 diode
R43717 N43716 N43717 10
D43717 N43717 0 diode
R43718 N43717 N43718 10
D43718 N43718 0 diode
R43719 N43718 N43719 10
D43719 N43719 0 diode
R43720 N43719 N43720 10
D43720 N43720 0 diode
R43721 N43720 N43721 10
D43721 N43721 0 diode
R43722 N43721 N43722 10
D43722 N43722 0 diode
R43723 N43722 N43723 10
D43723 N43723 0 diode
R43724 N43723 N43724 10
D43724 N43724 0 diode
R43725 N43724 N43725 10
D43725 N43725 0 diode
R43726 N43725 N43726 10
D43726 N43726 0 diode
R43727 N43726 N43727 10
D43727 N43727 0 diode
R43728 N43727 N43728 10
D43728 N43728 0 diode
R43729 N43728 N43729 10
D43729 N43729 0 diode
R43730 N43729 N43730 10
D43730 N43730 0 diode
R43731 N43730 N43731 10
D43731 N43731 0 diode
R43732 N43731 N43732 10
D43732 N43732 0 diode
R43733 N43732 N43733 10
D43733 N43733 0 diode
R43734 N43733 N43734 10
D43734 N43734 0 diode
R43735 N43734 N43735 10
D43735 N43735 0 diode
R43736 N43735 N43736 10
D43736 N43736 0 diode
R43737 N43736 N43737 10
D43737 N43737 0 diode
R43738 N43737 N43738 10
D43738 N43738 0 diode
R43739 N43738 N43739 10
D43739 N43739 0 diode
R43740 N43739 N43740 10
D43740 N43740 0 diode
R43741 N43740 N43741 10
D43741 N43741 0 diode
R43742 N43741 N43742 10
D43742 N43742 0 diode
R43743 N43742 N43743 10
D43743 N43743 0 diode
R43744 N43743 N43744 10
D43744 N43744 0 diode
R43745 N43744 N43745 10
D43745 N43745 0 diode
R43746 N43745 N43746 10
D43746 N43746 0 diode
R43747 N43746 N43747 10
D43747 N43747 0 diode
R43748 N43747 N43748 10
D43748 N43748 0 diode
R43749 N43748 N43749 10
D43749 N43749 0 diode
R43750 N43749 N43750 10
D43750 N43750 0 diode
R43751 N43750 N43751 10
D43751 N43751 0 diode
R43752 N43751 N43752 10
D43752 N43752 0 diode
R43753 N43752 N43753 10
D43753 N43753 0 diode
R43754 N43753 N43754 10
D43754 N43754 0 diode
R43755 N43754 N43755 10
D43755 N43755 0 diode
R43756 N43755 N43756 10
D43756 N43756 0 diode
R43757 N43756 N43757 10
D43757 N43757 0 diode
R43758 N43757 N43758 10
D43758 N43758 0 diode
R43759 N43758 N43759 10
D43759 N43759 0 diode
R43760 N43759 N43760 10
D43760 N43760 0 diode
R43761 N43760 N43761 10
D43761 N43761 0 diode
R43762 N43761 N43762 10
D43762 N43762 0 diode
R43763 N43762 N43763 10
D43763 N43763 0 diode
R43764 N43763 N43764 10
D43764 N43764 0 diode
R43765 N43764 N43765 10
D43765 N43765 0 diode
R43766 N43765 N43766 10
D43766 N43766 0 diode
R43767 N43766 N43767 10
D43767 N43767 0 diode
R43768 N43767 N43768 10
D43768 N43768 0 diode
R43769 N43768 N43769 10
D43769 N43769 0 diode
R43770 N43769 N43770 10
D43770 N43770 0 diode
R43771 N43770 N43771 10
D43771 N43771 0 diode
R43772 N43771 N43772 10
D43772 N43772 0 diode
R43773 N43772 N43773 10
D43773 N43773 0 diode
R43774 N43773 N43774 10
D43774 N43774 0 diode
R43775 N43774 N43775 10
D43775 N43775 0 diode
R43776 N43775 N43776 10
D43776 N43776 0 diode
R43777 N43776 N43777 10
D43777 N43777 0 diode
R43778 N43777 N43778 10
D43778 N43778 0 diode
R43779 N43778 N43779 10
D43779 N43779 0 diode
R43780 N43779 N43780 10
D43780 N43780 0 diode
R43781 N43780 N43781 10
D43781 N43781 0 diode
R43782 N43781 N43782 10
D43782 N43782 0 diode
R43783 N43782 N43783 10
D43783 N43783 0 diode
R43784 N43783 N43784 10
D43784 N43784 0 diode
R43785 N43784 N43785 10
D43785 N43785 0 diode
R43786 N43785 N43786 10
D43786 N43786 0 diode
R43787 N43786 N43787 10
D43787 N43787 0 diode
R43788 N43787 N43788 10
D43788 N43788 0 diode
R43789 N43788 N43789 10
D43789 N43789 0 diode
R43790 N43789 N43790 10
D43790 N43790 0 diode
R43791 N43790 N43791 10
D43791 N43791 0 diode
R43792 N43791 N43792 10
D43792 N43792 0 diode
R43793 N43792 N43793 10
D43793 N43793 0 diode
R43794 N43793 N43794 10
D43794 N43794 0 diode
R43795 N43794 N43795 10
D43795 N43795 0 diode
R43796 N43795 N43796 10
D43796 N43796 0 diode
R43797 N43796 N43797 10
D43797 N43797 0 diode
R43798 N43797 N43798 10
D43798 N43798 0 diode
R43799 N43798 N43799 10
D43799 N43799 0 diode
R43800 N43799 N43800 10
D43800 N43800 0 diode
R43801 N43800 N43801 10
D43801 N43801 0 diode
R43802 N43801 N43802 10
D43802 N43802 0 diode
R43803 N43802 N43803 10
D43803 N43803 0 diode
R43804 N43803 N43804 10
D43804 N43804 0 diode
R43805 N43804 N43805 10
D43805 N43805 0 diode
R43806 N43805 N43806 10
D43806 N43806 0 diode
R43807 N43806 N43807 10
D43807 N43807 0 diode
R43808 N43807 N43808 10
D43808 N43808 0 diode
R43809 N43808 N43809 10
D43809 N43809 0 diode
R43810 N43809 N43810 10
D43810 N43810 0 diode
R43811 N43810 N43811 10
D43811 N43811 0 diode
R43812 N43811 N43812 10
D43812 N43812 0 diode
R43813 N43812 N43813 10
D43813 N43813 0 diode
R43814 N43813 N43814 10
D43814 N43814 0 diode
R43815 N43814 N43815 10
D43815 N43815 0 diode
R43816 N43815 N43816 10
D43816 N43816 0 diode
R43817 N43816 N43817 10
D43817 N43817 0 diode
R43818 N43817 N43818 10
D43818 N43818 0 diode
R43819 N43818 N43819 10
D43819 N43819 0 diode
R43820 N43819 N43820 10
D43820 N43820 0 diode
R43821 N43820 N43821 10
D43821 N43821 0 diode
R43822 N43821 N43822 10
D43822 N43822 0 diode
R43823 N43822 N43823 10
D43823 N43823 0 diode
R43824 N43823 N43824 10
D43824 N43824 0 diode
R43825 N43824 N43825 10
D43825 N43825 0 diode
R43826 N43825 N43826 10
D43826 N43826 0 diode
R43827 N43826 N43827 10
D43827 N43827 0 diode
R43828 N43827 N43828 10
D43828 N43828 0 diode
R43829 N43828 N43829 10
D43829 N43829 0 diode
R43830 N43829 N43830 10
D43830 N43830 0 diode
R43831 N43830 N43831 10
D43831 N43831 0 diode
R43832 N43831 N43832 10
D43832 N43832 0 diode
R43833 N43832 N43833 10
D43833 N43833 0 diode
R43834 N43833 N43834 10
D43834 N43834 0 diode
R43835 N43834 N43835 10
D43835 N43835 0 diode
R43836 N43835 N43836 10
D43836 N43836 0 diode
R43837 N43836 N43837 10
D43837 N43837 0 diode
R43838 N43837 N43838 10
D43838 N43838 0 diode
R43839 N43838 N43839 10
D43839 N43839 0 diode
R43840 N43839 N43840 10
D43840 N43840 0 diode
R43841 N43840 N43841 10
D43841 N43841 0 diode
R43842 N43841 N43842 10
D43842 N43842 0 diode
R43843 N43842 N43843 10
D43843 N43843 0 diode
R43844 N43843 N43844 10
D43844 N43844 0 diode
R43845 N43844 N43845 10
D43845 N43845 0 diode
R43846 N43845 N43846 10
D43846 N43846 0 diode
R43847 N43846 N43847 10
D43847 N43847 0 diode
R43848 N43847 N43848 10
D43848 N43848 0 diode
R43849 N43848 N43849 10
D43849 N43849 0 diode
R43850 N43849 N43850 10
D43850 N43850 0 diode
R43851 N43850 N43851 10
D43851 N43851 0 diode
R43852 N43851 N43852 10
D43852 N43852 0 diode
R43853 N43852 N43853 10
D43853 N43853 0 diode
R43854 N43853 N43854 10
D43854 N43854 0 diode
R43855 N43854 N43855 10
D43855 N43855 0 diode
R43856 N43855 N43856 10
D43856 N43856 0 diode
R43857 N43856 N43857 10
D43857 N43857 0 diode
R43858 N43857 N43858 10
D43858 N43858 0 diode
R43859 N43858 N43859 10
D43859 N43859 0 diode
R43860 N43859 N43860 10
D43860 N43860 0 diode
R43861 N43860 N43861 10
D43861 N43861 0 diode
R43862 N43861 N43862 10
D43862 N43862 0 diode
R43863 N43862 N43863 10
D43863 N43863 0 diode
R43864 N43863 N43864 10
D43864 N43864 0 diode
R43865 N43864 N43865 10
D43865 N43865 0 diode
R43866 N43865 N43866 10
D43866 N43866 0 diode
R43867 N43866 N43867 10
D43867 N43867 0 diode
R43868 N43867 N43868 10
D43868 N43868 0 diode
R43869 N43868 N43869 10
D43869 N43869 0 diode
R43870 N43869 N43870 10
D43870 N43870 0 diode
R43871 N43870 N43871 10
D43871 N43871 0 diode
R43872 N43871 N43872 10
D43872 N43872 0 diode
R43873 N43872 N43873 10
D43873 N43873 0 diode
R43874 N43873 N43874 10
D43874 N43874 0 diode
R43875 N43874 N43875 10
D43875 N43875 0 diode
R43876 N43875 N43876 10
D43876 N43876 0 diode
R43877 N43876 N43877 10
D43877 N43877 0 diode
R43878 N43877 N43878 10
D43878 N43878 0 diode
R43879 N43878 N43879 10
D43879 N43879 0 diode
R43880 N43879 N43880 10
D43880 N43880 0 diode
R43881 N43880 N43881 10
D43881 N43881 0 diode
R43882 N43881 N43882 10
D43882 N43882 0 diode
R43883 N43882 N43883 10
D43883 N43883 0 diode
R43884 N43883 N43884 10
D43884 N43884 0 diode
R43885 N43884 N43885 10
D43885 N43885 0 diode
R43886 N43885 N43886 10
D43886 N43886 0 diode
R43887 N43886 N43887 10
D43887 N43887 0 diode
R43888 N43887 N43888 10
D43888 N43888 0 diode
R43889 N43888 N43889 10
D43889 N43889 0 diode
R43890 N43889 N43890 10
D43890 N43890 0 diode
R43891 N43890 N43891 10
D43891 N43891 0 diode
R43892 N43891 N43892 10
D43892 N43892 0 diode
R43893 N43892 N43893 10
D43893 N43893 0 diode
R43894 N43893 N43894 10
D43894 N43894 0 diode
R43895 N43894 N43895 10
D43895 N43895 0 diode
R43896 N43895 N43896 10
D43896 N43896 0 diode
R43897 N43896 N43897 10
D43897 N43897 0 diode
R43898 N43897 N43898 10
D43898 N43898 0 diode
R43899 N43898 N43899 10
D43899 N43899 0 diode
R43900 N43899 N43900 10
D43900 N43900 0 diode
R43901 N43900 N43901 10
D43901 N43901 0 diode
R43902 N43901 N43902 10
D43902 N43902 0 diode
R43903 N43902 N43903 10
D43903 N43903 0 diode
R43904 N43903 N43904 10
D43904 N43904 0 diode
R43905 N43904 N43905 10
D43905 N43905 0 diode
R43906 N43905 N43906 10
D43906 N43906 0 diode
R43907 N43906 N43907 10
D43907 N43907 0 diode
R43908 N43907 N43908 10
D43908 N43908 0 diode
R43909 N43908 N43909 10
D43909 N43909 0 diode
R43910 N43909 N43910 10
D43910 N43910 0 diode
R43911 N43910 N43911 10
D43911 N43911 0 diode
R43912 N43911 N43912 10
D43912 N43912 0 diode
R43913 N43912 N43913 10
D43913 N43913 0 diode
R43914 N43913 N43914 10
D43914 N43914 0 diode
R43915 N43914 N43915 10
D43915 N43915 0 diode
R43916 N43915 N43916 10
D43916 N43916 0 diode
R43917 N43916 N43917 10
D43917 N43917 0 diode
R43918 N43917 N43918 10
D43918 N43918 0 diode
R43919 N43918 N43919 10
D43919 N43919 0 diode
R43920 N43919 N43920 10
D43920 N43920 0 diode
R43921 N43920 N43921 10
D43921 N43921 0 diode
R43922 N43921 N43922 10
D43922 N43922 0 diode
R43923 N43922 N43923 10
D43923 N43923 0 diode
R43924 N43923 N43924 10
D43924 N43924 0 diode
R43925 N43924 N43925 10
D43925 N43925 0 diode
R43926 N43925 N43926 10
D43926 N43926 0 diode
R43927 N43926 N43927 10
D43927 N43927 0 diode
R43928 N43927 N43928 10
D43928 N43928 0 diode
R43929 N43928 N43929 10
D43929 N43929 0 diode
R43930 N43929 N43930 10
D43930 N43930 0 diode
R43931 N43930 N43931 10
D43931 N43931 0 diode
R43932 N43931 N43932 10
D43932 N43932 0 diode
R43933 N43932 N43933 10
D43933 N43933 0 diode
R43934 N43933 N43934 10
D43934 N43934 0 diode
R43935 N43934 N43935 10
D43935 N43935 0 diode
R43936 N43935 N43936 10
D43936 N43936 0 diode
R43937 N43936 N43937 10
D43937 N43937 0 diode
R43938 N43937 N43938 10
D43938 N43938 0 diode
R43939 N43938 N43939 10
D43939 N43939 0 diode
R43940 N43939 N43940 10
D43940 N43940 0 diode
R43941 N43940 N43941 10
D43941 N43941 0 diode
R43942 N43941 N43942 10
D43942 N43942 0 diode
R43943 N43942 N43943 10
D43943 N43943 0 diode
R43944 N43943 N43944 10
D43944 N43944 0 diode
R43945 N43944 N43945 10
D43945 N43945 0 diode
R43946 N43945 N43946 10
D43946 N43946 0 diode
R43947 N43946 N43947 10
D43947 N43947 0 diode
R43948 N43947 N43948 10
D43948 N43948 0 diode
R43949 N43948 N43949 10
D43949 N43949 0 diode
R43950 N43949 N43950 10
D43950 N43950 0 diode
R43951 N43950 N43951 10
D43951 N43951 0 diode
R43952 N43951 N43952 10
D43952 N43952 0 diode
R43953 N43952 N43953 10
D43953 N43953 0 diode
R43954 N43953 N43954 10
D43954 N43954 0 diode
R43955 N43954 N43955 10
D43955 N43955 0 diode
R43956 N43955 N43956 10
D43956 N43956 0 diode
R43957 N43956 N43957 10
D43957 N43957 0 diode
R43958 N43957 N43958 10
D43958 N43958 0 diode
R43959 N43958 N43959 10
D43959 N43959 0 diode
R43960 N43959 N43960 10
D43960 N43960 0 diode
R43961 N43960 N43961 10
D43961 N43961 0 diode
R43962 N43961 N43962 10
D43962 N43962 0 diode
R43963 N43962 N43963 10
D43963 N43963 0 diode
R43964 N43963 N43964 10
D43964 N43964 0 diode
R43965 N43964 N43965 10
D43965 N43965 0 diode
R43966 N43965 N43966 10
D43966 N43966 0 diode
R43967 N43966 N43967 10
D43967 N43967 0 diode
R43968 N43967 N43968 10
D43968 N43968 0 diode
R43969 N43968 N43969 10
D43969 N43969 0 diode
R43970 N43969 N43970 10
D43970 N43970 0 diode
R43971 N43970 N43971 10
D43971 N43971 0 diode
R43972 N43971 N43972 10
D43972 N43972 0 diode
R43973 N43972 N43973 10
D43973 N43973 0 diode
R43974 N43973 N43974 10
D43974 N43974 0 diode
R43975 N43974 N43975 10
D43975 N43975 0 diode
R43976 N43975 N43976 10
D43976 N43976 0 diode
R43977 N43976 N43977 10
D43977 N43977 0 diode
R43978 N43977 N43978 10
D43978 N43978 0 diode
R43979 N43978 N43979 10
D43979 N43979 0 diode
R43980 N43979 N43980 10
D43980 N43980 0 diode
R43981 N43980 N43981 10
D43981 N43981 0 diode
R43982 N43981 N43982 10
D43982 N43982 0 diode
R43983 N43982 N43983 10
D43983 N43983 0 diode
R43984 N43983 N43984 10
D43984 N43984 0 diode
R43985 N43984 N43985 10
D43985 N43985 0 diode
R43986 N43985 N43986 10
D43986 N43986 0 diode
R43987 N43986 N43987 10
D43987 N43987 0 diode
R43988 N43987 N43988 10
D43988 N43988 0 diode
R43989 N43988 N43989 10
D43989 N43989 0 diode
R43990 N43989 N43990 10
D43990 N43990 0 diode
R43991 N43990 N43991 10
D43991 N43991 0 diode
R43992 N43991 N43992 10
D43992 N43992 0 diode
R43993 N43992 N43993 10
D43993 N43993 0 diode
R43994 N43993 N43994 10
D43994 N43994 0 diode
R43995 N43994 N43995 10
D43995 N43995 0 diode
R43996 N43995 N43996 10
D43996 N43996 0 diode
R43997 N43996 N43997 10
D43997 N43997 0 diode
R43998 N43997 N43998 10
D43998 N43998 0 diode
R43999 N43998 N43999 10
D43999 N43999 0 diode
R44000 N43999 N44000 10
D44000 N44000 0 diode
R44001 N44000 N44001 10
D44001 N44001 0 diode
R44002 N44001 N44002 10
D44002 N44002 0 diode
R44003 N44002 N44003 10
D44003 N44003 0 diode
R44004 N44003 N44004 10
D44004 N44004 0 diode
R44005 N44004 N44005 10
D44005 N44005 0 diode
R44006 N44005 N44006 10
D44006 N44006 0 diode
R44007 N44006 N44007 10
D44007 N44007 0 diode
R44008 N44007 N44008 10
D44008 N44008 0 diode
R44009 N44008 N44009 10
D44009 N44009 0 diode
R44010 N44009 N44010 10
D44010 N44010 0 diode
R44011 N44010 N44011 10
D44011 N44011 0 diode
R44012 N44011 N44012 10
D44012 N44012 0 diode
R44013 N44012 N44013 10
D44013 N44013 0 diode
R44014 N44013 N44014 10
D44014 N44014 0 diode
R44015 N44014 N44015 10
D44015 N44015 0 diode
R44016 N44015 N44016 10
D44016 N44016 0 diode
R44017 N44016 N44017 10
D44017 N44017 0 diode
R44018 N44017 N44018 10
D44018 N44018 0 diode
R44019 N44018 N44019 10
D44019 N44019 0 diode
R44020 N44019 N44020 10
D44020 N44020 0 diode
R44021 N44020 N44021 10
D44021 N44021 0 diode
R44022 N44021 N44022 10
D44022 N44022 0 diode
R44023 N44022 N44023 10
D44023 N44023 0 diode
R44024 N44023 N44024 10
D44024 N44024 0 diode
R44025 N44024 N44025 10
D44025 N44025 0 diode
R44026 N44025 N44026 10
D44026 N44026 0 diode
R44027 N44026 N44027 10
D44027 N44027 0 diode
R44028 N44027 N44028 10
D44028 N44028 0 diode
R44029 N44028 N44029 10
D44029 N44029 0 diode
R44030 N44029 N44030 10
D44030 N44030 0 diode
R44031 N44030 N44031 10
D44031 N44031 0 diode
R44032 N44031 N44032 10
D44032 N44032 0 diode
R44033 N44032 N44033 10
D44033 N44033 0 diode
R44034 N44033 N44034 10
D44034 N44034 0 diode
R44035 N44034 N44035 10
D44035 N44035 0 diode
R44036 N44035 N44036 10
D44036 N44036 0 diode
R44037 N44036 N44037 10
D44037 N44037 0 diode
R44038 N44037 N44038 10
D44038 N44038 0 diode
R44039 N44038 N44039 10
D44039 N44039 0 diode
R44040 N44039 N44040 10
D44040 N44040 0 diode
R44041 N44040 N44041 10
D44041 N44041 0 diode
R44042 N44041 N44042 10
D44042 N44042 0 diode
R44043 N44042 N44043 10
D44043 N44043 0 diode
R44044 N44043 N44044 10
D44044 N44044 0 diode
R44045 N44044 N44045 10
D44045 N44045 0 diode
R44046 N44045 N44046 10
D44046 N44046 0 diode
R44047 N44046 N44047 10
D44047 N44047 0 diode
R44048 N44047 N44048 10
D44048 N44048 0 diode
R44049 N44048 N44049 10
D44049 N44049 0 diode
R44050 N44049 N44050 10
D44050 N44050 0 diode
R44051 N44050 N44051 10
D44051 N44051 0 diode
R44052 N44051 N44052 10
D44052 N44052 0 diode
R44053 N44052 N44053 10
D44053 N44053 0 diode
R44054 N44053 N44054 10
D44054 N44054 0 diode
R44055 N44054 N44055 10
D44055 N44055 0 diode
R44056 N44055 N44056 10
D44056 N44056 0 diode
R44057 N44056 N44057 10
D44057 N44057 0 diode
R44058 N44057 N44058 10
D44058 N44058 0 diode
R44059 N44058 N44059 10
D44059 N44059 0 diode
R44060 N44059 N44060 10
D44060 N44060 0 diode
R44061 N44060 N44061 10
D44061 N44061 0 diode
R44062 N44061 N44062 10
D44062 N44062 0 diode
R44063 N44062 N44063 10
D44063 N44063 0 diode
R44064 N44063 N44064 10
D44064 N44064 0 diode
R44065 N44064 N44065 10
D44065 N44065 0 diode
R44066 N44065 N44066 10
D44066 N44066 0 diode
R44067 N44066 N44067 10
D44067 N44067 0 diode
R44068 N44067 N44068 10
D44068 N44068 0 diode
R44069 N44068 N44069 10
D44069 N44069 0 diode
R44070 N44069 N44070 10
D44070 N44070 0 diode
R44071 N44070 N44071 10
D44071 N44071 0 diode
R44072 N44071 N44072 10
D44072 N44072 0 diode
R44073 N44072 N44073 10
D44073 N44073 0 diode
R44074 N44073 N44074 10
D44074 N44074 0 diode
R44075 N44074 N44075 10
D44075 N44075 0 diode
R44076 N44075 N44076 10
D44076 N44076 0 diode
R44077 N44076 N44077 10
D44077 N44077 0 diode
R44078 N44077 N44078 10
D44078 N44078 0 diode
R44079 N44078 N44079 10
D44079 N44079 0 diode
R44080 N44079 N44080 10
D44080 N44080 0 diode
R44081 N44080 N44081 10
D44081 N44081 0 diode
R44082 N44081 N44082 10
D44082 N44082 0 diode
R44083 N44082 N44083 10
D44083 N44083 0 diode
R44084 N44083 N44084 10
D44084 N44084 0 diode
R44085 N44084 N44085 10
D44085 N44085 0 diode
R44086 N44085 N44086 10
D44086 N44086 0 diode
R44087 N44086 N44087 10
D44087 N44087 0 diode
R44088 N44087 N44088 10
D44088 N44088 0 diode
R44089 N44088 N44089 10
D44089 N44089 0 diode
R44090 N44089 N44090 10
D44090 N44090 0 diode
R44091 N44090 N44091 10
D44091 N44091 0 diode
R44092 N44091 N44092 10
D44092 N44092 0 diode
R44093 N44092 N44093 10
D44093 N44093 0 diode
R44094 N44093 N44094 10
D44094 N44094 0 diode
R44095 N44094 N44095 10
D44095 N44095 0 diode
R44096 N44095 N44096 10
D44096 N44096 0 diode
R44097 N44096 N44097 10
D44097 N44097 0 diode
R44098 N44097 N44098 10
D44098 N44098 0 diode
R44099 N44098 N44099 10
D44099 N44099 0 diode
R44100 N44099 N44100 10
D44100 N44100 0 diode
R44101 N44100 N44101 10
D44101 N44101 0 diode
R44102 N44101 N44102 10
D44102 N44102 0 diode
R44103 N44102 N44103 10
D44103 N44103 0 diode
R44104 N44103 N44104 10
D44104 N44104 0 diode
R44105 N44104 N44105 10
D44105 N44105 0 diode
R44106 N44105 N44106 10
D44106 N44106 0 diode
R44107 N44106 N44107 10
D44107 N44107 0 diode
R44108 N44107 N44108 10
D44108 N44108 0 diode
R44109 N44108 N44109 10
D44109 N44109 0 diode
R44110 N44109 N44110 10
D44110 N44110 0 diode
R44111 N44110 N44111 10
D44111 N44111 0 diode
R44112 N44111 N44112 10
D44112 N44112 0 diode
R44113 N44112 N44113 10
D44113 N44113 0 diode
R44114 N44113 N44114 10
D44114 N44114 0 diode
R44115 N44114 N44115 10
D44115 N44115 0 diode
R44116 N44115 N44116 10
D44116 N44116 0 diode
R44117 N44116 N44117 10
D44117 N44117 0 diode
R44118 N44117 N44118 10
D44118 N44118 0 diode
R44119 N44118 N44119 10
D44119 N44119 0 diode
R44120 N44119 N44120 10
D44120 N44120 0 diode
R44121 N44120 N44121 10
D44121 N44121 0 diode
R44122 N44121 N44122 10
D44122 N44122 0 diode
R44123 N44122 N44123 10
D44123 N44123 0 diode
R44124 N44123 N44124 10
D44124 N44124 0 diode
R44125 N44124 N44125 10
D44125 N44125 0 diode
R44126 N44125 N44126 10
D44126 N44126 0 diode
R44127 N44126 N44127 10
D44127 N44127 0 diode
R44128 N44127 N44128 10
D44128 N44128 0 diode
R44129 N44128 N44129 10
D44129 N44129 0 diode
R44130 N44129 N44130 10
D44130 N44130 0 diode
R44131 N44130 N44131 10
D44131 N44131 0 diode
R44132 N44131 N44132 10
D44132 N44132 0 diode
R44133 N44132 N44133 10
D44133 N44133 0 diode
R44134 N44133 N44134 10
D44134 N44134 0 diode
R44135 N44134 N44135 10
D44135 N44135 0 diode
R44136 N44135 N44136 10
D44136 N44136 0 diode
R44137 N44136 N44137 10
D44137 N44137 0 diode
R44138 N44137 N44138 10
D44138 N44138 0 diode
R44139 N44138 N44139 10
D44139 N44139 0 diode
R44140 N44139 N44140 10
D44140 N44140 0 diode
R44141 N44140 N44141 10
D44141 N44141 0 diode
R44142 N44141 N44142 10
D44142 N44142 0 diode
R44143 N44142 N44143 10
D44143 N44143 0 diode
R44144 N44143 N44144 10
D44144 N44144 0 diode
R44145 N44144 N44145 10
D44145 N44145 0 diode
R44146 N44145 N44146 10
D44146 N44146 0 diode
R44147 N44146 N44147 10
D44147 N44147 0 diode
R44148 N44147 N44148 10
D44148 N44148 0 diode
R44149 N44148 N44149 10
D44149 N44149 0 diode
R44150 N44149 N44150 10
D44150 N44150 0 diode
R44151 N44150 N44151 10
D44151 N44151 0 diode
R44152 N44151 N44152 10
D44152 N44152 0 diode
R44153 N44152 N44153 10
D44153 N44153 0 diode
R44154 N44153 N44154 10
D44154 N44154 0 diode
R44155 N44154 N44155 10
D44155 N44155 0 diode
R44156 N44155 N44156 10
D44156 N44156 0 diode
R44157 N44156 N44157 10
D44157 N44157 0 diode
R44158 N44157 N44158 10
D44158 N44158 0 diode
R44159 N44158 N44159 10
D44159 N44159 0 diode
R44160 N44159 N44160 10
D44160 N44160 0 diode
R44161 N44160 N44161 10
D44161 N44161 0 diode
R44162 N44161 N44162 10
D44162 N44162 0 diode
R44163 N44162 N44163 10
D44163 N44163 0 diode
R44164 N44163 N44164 10
D44164 N44164 0 diode
R44165 N44164 N44165 10
D44165 N44165 0 diode
R44166 N44165 N44166 10
D44166 N44166 0 diode
R44167 N44166 N44167 10
D44167 N44167 0 diode
R44168 N44167 N44168 10
D44168 N44168 0 diode
R44169 N44168 N44169 10
D44169 N44169 0 diode
R44170 N44169 N44170 10
D44170 N44170 0 diode
R44171 N44170 N44171 10
D44171 N44171 0 diode
R44172 N44171 N44172 10
D44172 N44172 0 diode
R44173 N44172 N44173 10
D44173 N44173 0 diode
R44174 N44173 N44174 10
D44174 N44174 0 diode
R44175 N44174 N44175 10
D44175 N44175 0 diode
R44176 N44175 N44176 10
D44176 N44176 0 diode
R44177 N44176 N44177 10
D44177 N44177 0 diode
R44178 N44177 N44178 10
D44178 N44178 0 diode
R44179 N44178 N44179 10
D44179 N44179 0 diode
R44180 N44179 N44180 10
D44180 N44180 0 diode
R44181 N44180 N44181 10
D44181 N44181 0 diode
R44182 N44181 N44182 10
D44182 N44182 0 diode
R44183 N44182 N44183 10
D44183 N44183 0 diode
R44184 N44183 N44184 10
D44184 N44184 0 diode
R44185 N44184 N44185 10
D44185 N44185 0 diode
R44186 N44185 N44186 10
D44186 N44186 0 diode
R44187 N44186 N44187 10
D44187 N44187 0 diode
R44188 N44187 N44188 10
D44188 N44188 0 diode
R44189 N44188 N44189 10
D44189 N44189 0 diode
R44190 N44189 N44190 10
D44190 N44190 0 diode
R44191 N44190 N44191 10
D44191 N44191 0 diode
R44192 N44191 N44192 10
D44192 N44192 0 diode
R44193 N44192 N44193 10
D44193 N44193 0 diode
R44194 N44193 N44194 10
D44194 N44194 0 diode
R44195 N44194 N44195 10
D44195 N44195 0 diode
R44196 N44195 N44196 10
D44196 N44196 0 diode
R44197 N44196 N44197 10
D44197 N44197 0 diode
R44198 N44197 N44198 10
D44198 N44198 0 diode
R44199 N44198 N44199 10
D44199 N44199 0 diode
R44200 N44199 N44200 10
D44200 N44200 0 diode
R44201 N44200 N44201 10
D44201 N44201 0 diode
R44202 N44201 N44202 10
D44202 N44202 0 diode
R44203 N44202 N44203 10
D44203 N44203 0 diode
R44204 N44203 N44204 10
D44204 N44204 0 diode
R44205 N44204 N44205 10
D44205 N44205 0 diode
R44206 N44205 N44206 10
D44206 N44206 0 diode
R44207 N44206 N44207 10
D44207 N44207 0 diode
R44208 N44207 N44208 10
D44208 N44208 0 diode
R44209 N44208 N44209 10
D44209 N44209 0 diode
R44210 N44209 N44210 10
D44210 N44210 0 diode
R44211 N44210 N44211 10
D44211 N44211 0 diode
R44212 N44211 N44212 10
D44212 N44212 0 diode
R44213 N44212 N44213 10
D44213 N44213 0 diode
R44214 N44213 N44214 10
D44214 N44214 0 diode
R44215 N44214 N44215 10
D44215 N44215 0 diode
R44216 N44215 N44216 10
D44216 N44216 0 diode
R44217 N44216 N44217 10
D44217 N44217 0 diode
R44218 N44217 N44218 10
D44218 N44218 0 diode
R44219 N44218 N44219 10
D44219 N44219 0 diode
R44220 N44219 N44220 10
D44220 N44220 0 diode
R44221 N44220 N44221 10
D44221 N44221 0 diode
R44222 N44221 N44222 10
D44222 N44222 0 diode
R44223 N44222 N44223 10
D44223 N44223 0 diode
R44224 N44223 N44224 10
D44224 N44224 0 diode
R44225 N44224 N44225 10
D44225 N44225 0 diode
R44226 N44225 N44226 10
D44226 N44226 0 diode
R44227 N44226 N44227 10
D44227 N44227 0 diode
R44228 N44227 N44228 10
D44228 N44228 0 diode
R44229 N44228 N44229 10
D44229 N44229 0 diode
R44230 N44229 N44230 10
D44230 N44230 0 diode
R44231 N44230 N44231 10
D44231 N44231 0 diode
R44232 N44231 N44232 10
D44232 N44232 0 diode
R44233 N44232 N44233 10
D44233 N44233 0 diode
R44234 N44233 N44234 10
D44234 N44234 0 diode
R44235 N44234 N44235 10
D44235 N44235 0 diode
R44236 N44235 N44236 10
D44236 N44236 0 diode
R44237 N44236 N44237 10
D44237 N44237 0 diode
R44238 N44237 N44238 10
D44238 N44238 0 diode
R44239 N44238 N44239 10
D44239 N44239 0 diode
R44240 N44239 N44240 10
D44240 N44240 0 diode
R44241 N44240 N44241 10
D44241 N44241 0 diode
R44242 N44241 N44242 10
D44242 N44242 0 diode
R44243 N44242 N44243 10
D44243 N44243 0 diode
R44244 N44243 N44244 10
D44244 N44244 0 diode
R44245 N44244 N44245 10
D44245 N44245 0 diode
R44246 N44245 N44246 10
D44246 N44246 0 diode
R44247 N44246 N44247 10
D44247 N44247 0 diode
R44248 N44247 N44248 10
D44248 N44248 0 diode
R44249 N44248 N44249 10
D44249 N44249 0 diode
R44250 N44249 N44250 10
D44250 N44250 0 diode
R44251 N44250 N44251 10
D44251 N44251 0 diode
R44252 N44251 N44252 10
D44252 N44252 0 diode
R44253 N44252 N44253 10
D44253 N44253 0 diode
R44254 N44253 N44254 10
D44254 N44254 0 diode
R44255 N44254 N44255 10
D44255 N44255 0 diode
R44256 N44255 N44256 10
D44256 N44256 0 diode
R44257 N44256 N44257 10
D44257 N44257 0 diode
R44258 N44257 N44258 10
D44258 N44258 0 diode
R44259 N44258 N44259 10
D44259 N44259 0 diode
R44260 N44259 N44260 10
D44260 N44260 0 diode
R44261 N44260 N44261 10
D44261 N44261 0 diode
R44262 N44261 N44262 10
D44262 N44262 0 diode
R44263 N44262 N44263 10
D44263 N44263 0 diode
R44264 N44263 N44264 10
D44264 N44264 0 diode
R44265 N44264 N44265 10
D44265 N44265 0 diode
R44266 N44265 N44266 10
D44266 N44266 0 diode
R44267 N44266 N44267 10
D44267 N44267 0 diode
R44268 N44267 N44268 10
D44268 N44268 0 diode
R44269 N44268 N44269 10
D44269 N44269 0 diode
R44270 N44269 N44270 10
D44270 N44270 0 diode
R44271 N44270 N44271 10
D44271 N44271 0 diode
R44272 N44271 N44272 10
D44272 N44272 0 diode
R44273 N44272 N44273 10
D44273 N44273 0 diode
R44274 N44273 N44274 10
D44274 N44274 0 diode
R44275 N44274 N44275 10
D44275 N44275 0 diode
R44276 N44275 N44276 10
D44276 N44276 0 diode
R44277 N44276 N44277 10
D44277 N44277 0 diode
R44278 N44277 N44278 10
D44278 N44278 0 diode
R44279 N44278 N44279 10
D44279 N44279 0 diode
R44280 N44279 N44280 10
D44280 N44280 0 diode
R44281 N44280 N44281 10
D44281 N44281 0 diode
R44282 N44281 N44282 10
D44282 N44282 0 diode
R44283 N44282 N44283 10
D44283 N44283 0 diode
R44284 N44283 N44284 10
D44284 N44284 0 diode
R44285 N44284 N44285 10
D44285 N44285 0 diode
R44286 N44285 N44286 10
D44286 N44286 0 diode
R44287 N44286 N44287 10
D44287 N44287 0 diode
R44288 N44287 N44288 10
D44288 N44288 0 diode
R44289 N44288 N44289 10
D44289 N44289 0 diode
R44290 N44289 N44290 10
D44290 N44290 0 diode
R44291 N44290 N44291 10
D44291 N44291 0 diode
R44292 N44291 N44292 10
D44292 N44292 0 diode
R44293 N44292 N44293 10
D44293 N44293 0 diode
R44294 N44293 N44294 10
D44294 N44294 0 diode
R44295 N44294 N44295 10
D44295 N44295 0 diode
R44296 N44295 N44296 10
D44296 N44296 0 diode
R44297 N44296 N44297 10
D44297 N44297 0 diode
R44298 N44297 N44298 10
D44298 N44298 0 diode
R44299 N44298 N44299 10
D44299 N44299 0 diode
R44300 N44299 N44300 10
D44300 N44300 0 diode
R44301 N44300 N44301 10
D44301 N44301 0 diode
R44302 N44301 N44302 10
D44302 N44302 0 diode
R44303 N44302 N44303 10
D44303 N44303 0 diode
R44304 N44303 N44304 10
D44304 N44304 0 diode
R44305 N44304 N44305 10
D44305 N44305 0 diode
R44306 N44305 N44306 10
D44306 N44306 0 diode
R44307 N44306 N44307 10
D44307 N44307 0 diode
R44308 N44307 N44308 10
D44308 N44308 0 diode
R44309 N44308 N44309 10
D44309 N44309 0 diode
R44310 N44309 N44310 10
D44310 N44310 0 diode
R44311 N44310 N44311 10
D44311 N44311 0 diode
R44312 N44311 N44312 10
D44312 N44312 0 diode
R44313 N44312 N44313 10
D44313 N44313 0 diode
R44314 N44313 N44314 10
D44314 N44314 0 diode
R44315 N44314 N44315 10
D44315 N44315 0 diode
R44316 N44315 N44316 10
D44316 N44316 0 diode
R44317 N44316 N44317 10
D44317 N44317 0 diode
R44318 N44317 N44318 10
D44318 N44318 0 diode
R44319 N44318 N44319 10
D44319 N44319 0 diode
R44320 N44319 N44320 10
D44320 N44320 0 diode
R44321 N44320 N44321 10
D44321 N44321 0 diode
R44322 N44321 N44322 10
D44322 N44322 0 diode
R44323 N44322 N44323 10
D44323 N44323 0 diode
R44324 N44323 N44324 10
D44324 N44324 0 diode
R44325 N44324 N44325 10
D44325 N44325 0 diode
R44326 N44325 N44326 10
D44326 N44326 0 diode
R44327 N44326 N44327 10
D44327 N44327 0 diode
R44328 N44327 N44328 10
D44328 N44328 0 diode
R44329 N44328 N44329 10
D44329 N44329 0 diode
R44330 N44329 N44330 10
D44330 N44330 0 diode
R44331 N44330 N44331 10
D44331 N44331 0 diode
R44332 N44331 N44332 10
D44332 N44332 0 diode
R44333 N44332 N44333 10
D44333 N44333 0 diode
R44334 N44333 N44334 10
D44334 N44334 0 diode
R44335 N44334 N44335 10
D44335 N44335 0 diode
R44336 N44335 N44336 10
D44336 N44336 0 diode
R44337 N44336 N44337 10
D44337 N44337 0 diode
R44338 N44337 N44338 10
D44338 N44338 0 diode
R44339 N44338 N44339 10
D44339 N44339 0 diode
R44340 N44339 N44340 10
D44340 N44340 0 diode
R44341 N44340 N44341 10
D44341 N44341 0 diode
R44342 N44341 N44342 10
D44342 N44342 0 diode
R44343 N44342 N44343 10
D44343 N44343 0 diode
R44344 N44343 N44344 10
D44344 N44344 0 diode
R44345 N44344 N44345 10
D44345 N44345 0 diode
R44346 N44345 N44346 10
D44346 N44346 0 diode
R44347 N44346 N44347 10
D44347 N44347 0 diode
R44348 N44347 N44348 10
D44348 N44348 0 diode
R44349 N44348 N44349 10
D44349 N44349 0 diode
R44350 N44349 N44350 10
D44350 N44350 0 diode
R44351 N44350 N44351 10
D44351 N44351 0 diode
R44352 N44351 N44352 10
D44352 N44352 0 diode
R44353 N44352 N44353 10
D44353 N44353 0 diode
R44354 N44353 N44354 10
D44354 N44354 0 diode
R44355 N44354 N44355 10
D44355 N44355 0 diode
R44356 N44355 N44356 10
D44356 N44356 0 diode
R44357 N44356 N44357 10
D44357 N44357 0 diode
R44358 N44357 N44358 10
D44358 N44358 0 diode
R44359 N44358 N44359 10
D44359 N44359 0 diode
R44360 N44359 N44360 10
D44360 N44360 0 diode
R44361 N44360 N44361 10
D44361 N44361 0 diode
R44362 N44361 N44362 10
D44362 N44362 0 diode
R44363 N44362 N44363 10
D44363 N44363 0 diode
R44364 N44363 N44364 10
D44364 N44364 0 diode
R44365 N44364 N44365 10
D44365 N44365 0 diode
R44366 N44365 N44366 10
D44366 N44366 0 diode
R44367 N44366 N44367 10
D44367 N44367 0 diode
R44368 N44367 N44368 10
D44368 N44368 0 diode
R44369 N44368 N44369 10
D44369 N44369 0 diode
R44370 N44369 N44370 10
D44370 N44370 0 diode
R44371 N44370 N44371 10
D44371 N44371 0 diode
R44372 N44371 N44372 10
D44372 N44372 0 diode
R44373 N44372 N44373 10
D44373 N44373 0 diode
R44374 N44373 N44374 10
D44374 N44374 0 diode
R44375 N44374 N44375 10
D44375 N44375 0 diode
R44376 N44375 N44376 10
D44376 N44376 0 diode
R44377 N44376 N44377 10
D44377 N44377 0 diode
R44378 N44377 N44378 10
D44378 N44378 0 diode
R44379 N44378 N44379 10
D44379 N44379 0 diode
R44380 N44379 N44380 10
D44380 N44380 0 diode
R44381 N44380 N44381 10
D44381 N44381 0 diode
R44382 N44381 N44382 10
D44382 N44382 0 diode
R44383 N44382 N44383 10
D44383 N44383 0 diode
R44384 N44383 N44384 10
D44384 N44384 0 diode
R44385 N44384 N44385 10
D44385 N44385 0 diode
R44386 N44385 N44386 10
D44386 N44386 0 diode
R44387 N44386 N44387 10
D44387 N44387 0 diode
R44388 N44387 N44388 10
D44388 N44388 0 diode
R44389 N44388 N44389 10
D44389 N44389 0 diode
R44390 N44389 N44390 10
D44390 N44390 0 diode
R44391 N44390 N44391 10
D44391 N44391 0 diode
R44392 N44391 N44392 10
D44392 N44392 0 diode
R44393 N44392 N44393 10
D44393 N44393 0 diode
R44394 N44393 N44394 10
D44394 N44394 0 diode
R44395 N44394 N44395 10
D44395 N44395 0 diode
R44396 N44395 N44396 10
D44396 N44396 0 diode
R44397 N44396 N44397 10
D44397 N44397 0 diode
R44398 N44397 N44398 10
D44398 N44398 0 diode
R44399 N44398 N44399 10
D44399 N44399 0 diode
R44400 N44399 N44400 10
D44400 N44400 0 diode
R44401 N44400 N44401 10
D44401 N44401 0 diode
R44402 N44401 N44402 10
D44402 N44402 0 diode
R44403 N44402 N44403 10
D44403 N44403 0 diode
R44404 N44403 N44404 10
D44404 N44404 0 diode
R44405 N44404 N44405 10
D44405 N44405 0 diode
R44406 N44405 N44406 10
D44406 N44406 0 diode
R44407 N44406 N44407 10
D44407 N44407 0 diode
R44408 N44407 N44408 10
D44408 N44408 0 diode
R44409 N44408 N44409 10
D44409 N44409 0 diode
R44410 N44409 N44410 10
D44410 N44410 0 diode
R44411 N44410 N44411 10
D44411 N44411 0 diode
R44412 N44411 N44412 10
D44412 N44412 0 diode
R44413 N44412 N44413 10
D44413 N44413 0 diode
R44414 N44413 N44414 10
D44414 N44414 0 diode
R44415 N44414 N44415 10
D44415 N44415 0 diode
R44416 N44415 N44416 10
D44416 N44416 0 diode
R44417 N44416 N44417 10
D44417 N44417 0 diode
R44418 N44417 N44418 10
D44418 N44418 0 diode
R44419 N44418 N44419 10
D44419 N44419 0 diode
R44420 N44419 N44420 10
D44420 N44420 0 diode
R44421 N44420 N44421 10
D44421 N44421 0 diode
R44422 N44421 N44422 10
D44422 N44422 0 diode
R44423 N44422 N44423 10
D44423 N44423 0 diode
R44424 N44423 N44424 10
D44424 N44424 0 diode
R44425 N44424 N44425 10
D44425 N44425 0 diode
R44426 N44425 N44426 10
D44426 N44426 0 diode
R44427 N44426 N44427 10
D44427 N44427 0 diode
R44428 N44427 N44428 10
D44428 N44428 0 diode
R44429 N44428 N44429 10
D44429 N44429 0 diode
R44430 N44429 N44430 10
D44430 N44430 0 diode
R44431 N44430 N44431 10
D44431 N44431 0 diode
R44432 N44431 N44432 10
D44432 N44432 0 diode
R44433 N44432 N44433 10
D44433 N44433 0 diode
R44434 N44433 N44434 10
D44434 N44434 0 diode
R44435 N44434 N44435 10
D44435 N44435 0 diode
R44436 N44435 N44436 10
D44436 N44436 0 diode
R44437 N44436 N44437 10
D44437 N44437 0 diode
R44438 N44437 N44438 10
D44438 N44438 0 diode
R44439 N44438 N44439 10
D44439 N44439 0 diode
R44440 N44439 N44440 10
D44440 N44440 0 diode
R44441 N44440 N44441 10
D44441 N44441 0 diode
R44442 N44441 N44442 10
D44442 N44442 0 diode
R44443 N44442 N44443 10
D44443 N44443 0 diode
R44444 N44443 N44444 10
D44444 N44444 0 diode
R44445 N44444 N44445 10
D44445 N44445 0 diode
R44446 N44445 N44446 10
D44446 N44446 0 diode
R44447 N44446 N44447 10
D44447 N44447 0 diode
R44448 N44447 N44448 10
D44448 N44448 0 diode
R44449 N44448 N44449 10
D44449 N44449 0 diode
R44450 N44449 N44450 10
D44450 N44450 0 diode
R44451 N44450 N44451 10
D44451 N44451 0 diode
R44452 N44451 N44452 10
D44452 N44452 0 diode
R44453 N44452 N44453 10
D44453 N44453 0 diode
R44454 N44453 N44454 10
D44454 N44454 0 diode
R44455 N44454 N44455 10
D44455 N44455 0 diode
R44456 N44455 N44456 10
D44456 N44456 0 diode
R44457 N44456 N44457 10
D44457 N44457 0 diode
R44458 N44457 N44458 10
D44458 N44458 0 diode
R44459 N44458 N44459 10
D44459 N44459 0 diode
R44460 N44459 N44460 10
D44460 N44460 0 diode
R44461 N44460 N44461 10
D44461 N44461 0 diode
R44462 N44461 N44462 10
D44462 N44462 0 diode
R44463 N44462 N44463 10
D44463 N44463 0 diode
R44464 N44463 N44464 10
D44464 N44464 0 diode
R44465 N44464 N44465 10
D44465 N44465 0 diode
R44466 N44465 N44466 10
D44466 N44466 0 diode
R44467 N44466 N44467 10
D44467 N44467 0 diode
R44468 N44467 N44468 10
D44468 N44468 0 diode
R44469 N44468 N44469 10
D44469 N44469 0 diode
R44470 N44469 N44470 10
D44470 N44470 0 diode
R44471 N44470 N44471 10
D44471 N44471 0 diode
R44472 N44471 N44472 10
D44472 N44472 0 diode
R44473 N44472 N44473 10
D44473 N44473 0 diode
R44474 N44473 N44474 10
D44474 N44474 0 diode
R44475 N44474 N44475 10
D44475 N44475 0 diode
R44476 N44475 N44476 10
D44476 N44476 0 diode
R44477 N44476 N44477 10
D44477 N44477 0 diode
R44478 N44477 N44478 10
D44478 N44478 0 diode
R44479 N44478 N44479 10
D44479 N44479 0 diode
R44480 N44479 N44480 10
D44480 N44480 0 diode
R44481 N44480 N44481 10
D44481 N44481 0 diode
R44482 N44481 N44482 10
D44482 N44482 0 diode
R44483 N44482 N44483 10
D44483 N44483 0 diode
R44484 N44483 N44484 10
D44484 N44484 0 diode
R44485 N44484 N44485 10
D44485 N44485 0 diode
R44486 N44485 N44486 10
D44486 N44486 0 diode
R44487 N44486 N44487 10
D44487 N44487 0 diode
R44488 N44487 N44488 10
D44488 N44488 0 diode
R44489 N44488 N44489 10
D44489 N44489 0 diode
R44490 N44489 N44490 10
D44490 N44490 0 diode
R44491 N44490 N44491 10
D44491 N44491 0 diode
R44492 N44491 N44492 10
D44492 N44492 0 diode
R44493 N44492 N44493 10
D44493 N44493 0 diode
R44494 N44493 N44494 10
D44494 N44494 0 diode
R44495 N44494 N44495 10
D44495 N44495 0 diode
R44496 N44495 N44496 10
D44496 N44496 0 diode
R44497 N44496 N44497 10
D44497 N44497 0 diode
R44498 N44497 N44498 10
D44498 N44498 0 diode
R44499 N44498 N44499 10
D44499 N44499 0 diode
R44500 N44499 N44500 10
D44500 N44500 0 diode
R44501 N44500 N44501 10
D44501 N44501 0 diode
R44502 N44501 N44502 10
D44502 N44502 0 diode
R44503 N44502 N44503 10
D44503 N44503 0 diode
R44504 N44503 N44504 10
D44504 N44504 0 diode
R44505 N44504 N44505 10
D44505 N44505 0 diode
R44506 N44505 N44506 10
D44506 N44506 0 diode
R44507 N44506 N44507 10
D44507 N44507 0 diode
R44508 N44507 N44508 10
D44508 N44508 0 diode
R44509 N44508 N44509 10
D44509 N44509 0 diode
R44510 N44509 N44510 10
D44510 N44510 0 diode
R44511 N44510 N44511 10
D44511 N44511 0 diode
R44512 N44511 N44512 10
D44512 N44512 0 diode
R44513 N44512 N44513 10
D44513 N44513 0 diode
R44514 N44513 N44514 10
D44514 N44514 0 diode
R44515 N44514 N44515 10
D44515 N44515 0 diode
R44516 N44515 N44516 10
D44516 N44516 0 diode
R44517 N44516 N44517 10
D44517 N44517 0 diode
R44518 N44517 N44518 10
D44518 N44518 0 diode
R44519 N44518 N44519 10
D44519 N44519 0 diode
R44520 N44519 N44520 10
D44520 N44520 0 diode
R44521 N44520 N44521 10
D44521 N44521 0 diode
R44522 N44521 N44522 10
D44522 N44522 0 diode
R44523 N44522 N44523 10
D44523 N44523 0 diode
R44524 N44523 N44524 10
D44524 N44524 0 diode
R44525 N44524 N44525 10
D44525 N44525 0 diode
R44526 N44525 N44526 10
D44526 N44526 0 diode
R44527 N44526 N44527 10
D44527 N44527 0 diode
R44528 N44527 N44528 10
D44528 N44528 0 diode
R44529 N44528 N44529 10
D44529 N44529 0 diode
R44530 N44529 N44530 10
D44530 N44530 0 diode
R44531 N44530 N44531 10
D44531 N44531 0 diode
R44532 N44531 N44532 10
D44532 N44532 0 diode
R44533 N44532 N44533 10
D44533 N44533 0 diode
R44534 N44533 N44534 10
D44534 N44534 0 diode
R44535 N44534 N44535 10
D44535 N44535 0 diode
R44536 N44535 N44536 10
D44536 N44536 0 diode
R44537 N44536 N44537 10
D44537 N44537 0 diode
R44538 N44537 N44538 10
D44538 N44538 0 diode
R44539 N44538 N44539 10
D44539 N44539 0 diode
R44540 N44539 N44540 10
D44540 N44540 0 diode
R44541 N44540 N44541 10
D44541 N44541 0 diode
R44542 N44541 N44542 10
D44542 N44542 0 diode
R44543 N44542 N44543 10
D44543 N44543 0 diode
R44544 N44543 N44544 10
D44544 N44544 0 diode
R44545 N44544 N44545 10
D44545 N44545 0 diode
R44546 N44545 N44546 10
D44546 N44546 0 diode
R44547 N44546 N44547 10
D44547 N44547 0 diode
R44548 N44547 N44548 10
D44548 N44548 0 diode
R44549 N44548 N44549 10
D44549 N44549 0 diode
R44550 N44549 N44550 10
D44550 N44550 0 diode
R44551 N44550 N44551 10
D44551 N44551 0 diode
R44552 N44551 N44552 10
D44552 N44552 0 diode
R44553 N44552 N44553 10
D44553 N44553 0 diode
R44554 N44553 N44554 10
D44554 N44554 0 diode
R44555 N44554 N44555 10
D44555 N44555 0 diode
R44556 N44555 N44556 10
D44556 N44556 0 diode
R44557 N44556 N44557 10
D44557 N44557 0 diode
R44558 N44557 N44558 10
D44558 N44558 0 diode
R44559 N44558 N44559 10
D44559 N44559 0 diode
R44560 N44559 N44560 10
D44560 N44560 0 diode
R44561 N44560 N44561 10
D44561 N44561 0 diode
R44562 N44561 N44562 10
D44562 N44562 0 diode
R44563 N44562 N44563 10
D44563 N44563 0 diode
R44564 N44563 N44564 10
D44564 N44564 0 diode
R44565 N44564 N44565 10
D44565 N44565 0 diode
R44566 N44565 N44566 10
D44566 N44566 0 diode
R44567 N44566 N44567 10
D44567 N44567 0 diode
R44568 N44567 N44568 10
D44568 N44568 0 diode
R44569 N44568 N44569 10
D44569 N44569 0 diode
R44570 N44569 N44570 10
D44570 N44570 0 diode
R44571 N44570 N44571 10
D44571 N44571 0 diode
R44572 N44571 N44572 10
D44572 N44572 0 diode
R44573 N44572 N44573 10
D44573 N44573 0 diode
R44574 N44573 N44574 10
D44574 N44574 0 diode
R44575 N44574 N44575 10
D44575 N44575 0 diode
R44576 N44575 N44576 10
D44576 N44576 0 diode
R44577 N44576 N44577 10
D44577 N44577 0 diode
R44578 N44577 N44578 10
D44578 N44578 0 diode
R44579 N44578 N44579 10
D44579 N44579 0 diode
R44580 N44579 N44580 10
D44580 N44580 0 diode
R44581 N44580 N44581 10
D44581 N44581 0 diode
R44582 N44581 N44582 10
D44582 N44582 0 diode
R44583 N44582 N44583 10
D44583 N44583 0 diode
R44584 N44583 N44584 10
D44584 N44584 0 diode
R44585 N44584 N44585 10
D44585 N44585 0 diode
R44586 N44585 N44586 10
D44586 N44586 0 diode
R44587 N44586 N44587 10
D44587 N44587 0 diode
R44588 N44587 N44588 10
D44588 N44588 0 diode
R44589 N44588 N44589 10
D44589 N44589 0 diode
R44590 N44589 N44590 10
D44590 N44590 0 diode
R44591 N44590 N44591 10
D44591 N44591 0 diode
R44592 N44591 N44592 10
D44592 N44592 0 diode
R44593 N44592 N44593 10
D44593 N44593 0 diode
R44594 N44593 N44594 10
D44594 N44594 0 diode
R44595 N44594 N44595 10
D44595 N44595 0 diode
R44596 N44595 N44596 10
D44596 N44596 0 diode
R44597 N44596 N44597 10
D44597 N44597 0 diode
R44598 N44597 N44598 10
D44598 N44598 0 diode
R44599 N44598 N44599 10
D44599 N44599 0 diode
R44600 N44599 N44600 10
D44600 N44600 0 diode
R44601 N44600 N44601 10
D44601 N44601 0 diode
R44602 N44601 N44602 10
D44602 N44602 0 diode
R44603 N44602 N44603 10
D44603 N44603 0 diode
R44604 N44603 N44604 10
D44604 N44604 0 diode
R44605 N44604 N44605 10
D44605 N44605 0 diode
R44606 N44605 N44606 10
D44606 N44606 0 diode
R44607 N44606 N44607 10
D44607 N44607 0 diode
R44608 N44607 N44608 10
D44608 N44608 0 diode
R44609 N44608 N44609 10
D44609 N44609 0 diode
R44610 N44609 N44610 10
D44610 N44610 0 diode
R44611 N44610 N44611 10
D44611 N44611 0 diode
R44612 N44611 N44612 10
D44612 N44612 0 diode
R44613 N44612 N44613 10
D44613 N44613 0 diode
R44614 N44613 N44614 10
D44614 N44614 0 diode
R44615 N44614 N44615 10
D44615 N44615 0 diode
R44616 N44615 N44616 10
D44616 N44616 0 diode
R44617 N44616 N44617 10
D44617 N44617 0 diode
R44618 N44617 N44618 10
D44618 N44618 0 diode
R44619 N44618 N44619 10
D44619 N44619 0 diode
R44620 N44619 N44620 10
D44620 N44620 0 diode
R44621 N44620 N44621 10
D44621 N44621 0 diode
R44622 N44621 N44622 10
D44622 N44622 0 diode
R44623 N44622 N44623 10
D44623 N44623 0 diode
R44624 N44623 N44624 10
D44624 N44624 0 diode
R44625 N44624 N44625 10
D44625 N44625 0 diode
R44626 N44625 N44626 10
D44626 N44626 0 diode
R44627 N44626 N44627 10
D44627 N44627 0 diode
R44628 N44627 N44628 10
D44628 N44628 0 diode
R44629 N44628 N44629 10
D44629 N44629 0 diode
R44630 N44629 N44630 10
D44630 N44630 0 diode
R44631 N44630 N44631 10
D44631 N44631 0 diode
R44632 N44631 N44632 10
D44632 N44632 0 diode
R44633 N44632 N44633 10
D44633 N44633 0 diode
R44634 N44633 N44634 10
D44634 N44634 0 diode
R44635 N44634 N44635 10
D44635 N44635 0 diode
R44636 N44635 N44636 10
D44636 N44636 0 diode
R44637 N44636 N44637 10
D44637 N44637 0 diode
R44638 N44637 N44638 10
D44638 N44638 0 diode
R44639 N44638 N44639 10
D44639 N44639 0 diode
R44640 N44639 N44640 10
D44640 N44640 0 diode
R44641 N44640 N44641 10
D44641 N44641 0 diode
R44642 N44641 N44642 10
D44642 N44642 0 diode
R44643 N44642 N44643 10
D44643 N44643 0 diode
R44644 N44643 N44644 10
D44644 N44644 0 diode
R44645 N44644 N44645 10
D44645 N44645 0 diode
R44646 N44645 N44646 10
D44646 N44646 0 diode
R44647 N44646 N44647 10
D44647 N44647 0 diode
R44648 N44647 N44648 10
D44648 N44648 0 diode
R44649 N44648 N44649 10
D44649 N44649 0 diode
R44650 N44649 N44650 10
D44650 N44650 0 diode
R44651 N44650 N44651 10
D44651 N44651 0 diode
R44652 N44651 N44652 10
D44652 N44652 0 diode
R44653 N44652 N44653 10
D44653 N44653 0 diode
R44654 N44653 N44654 10
D44654 N44654 0 diode
R44655 N44654 N44655 10
D44655 N44655 0 diode
R44656 N44655 N44656 10
D44656 N44656 0 diode
R44657 N44656 N44657 10
D44657 N44657 0 diode
R44658 N44657 N44658 10
D44658 N44658 0 diode
R44659 N44658 N44659 10
D44659 N44659 0 diode
R44660 N44659 N44660 10
D44660 N44660 0 diode
R44661 N44660 N44661 10
D44661 N44661 0 diode
R44662 N44661 N44662 10
D44662 N44662 0 diode
R44663 N44662 N44663 10
D44663 N44663 0 diode
R44664 N44663 N44664 10
D44664 N44664 0 diode
R44665 N44664 N44665 10
D44665 N44665 0 diode
R44666 N44665 N44666 10
D44666 N44666 0 diode
R44667 N44666 N44667 10
D44667 N44667 0 diode
R44668 N44667 N44668 10
D44668 N44668 0 diode
R44669 N44668 N44669 10
D44669 N44669 0 diode
R44670 N44669 N44670 10
D44670 N44670 0 diode
R44671 N44670 N44671 10
D44671 N44671 0 diode
R44672 N44671 N44672 10
D44672 N44672 0 diode
R44673 N44672 N44673 10
D44673 N44673 0 diode
R44674 N44673 N44674 10
D44674 N44674 0 diode
R44675 N44674 N44675 10
D44675 N44675 0 diode
R44676 N44675 N44676 10
D44676 N44676 0 diode
R44677 N44676 N44677 10
D44677 N44677 0 diode
R44678 N44677 N44678 10
D44678 N44678 0 diode
R44679 N44678 N44679 10
D44679 N44679 0 diode
R44680 N44679 N44680 10
D44680 N44680 0 diode
R44681 N44680 N44681 10
D44681 N44681 0 diode
R44682 N44681 N44682 10
D44682 N44682 0 diode
R44683 N44682 N44683 10
D44683 N44683 0 diode
R44684 N44683 N44684 10
D44684 N44684 0 diode
R44685 N44684 N44685 10
D44685 N44685 0 diode
R44686 N44685 N44686 10
D44686 N44686 0 diode
R44687 N44686 N44687 10
D44687 N44687 0 diode
R44688 N44687 N44688 10
D44688 N44688 0 diode
R44689 N44688 N44689 10
D44689 N44689 0 diode
R44690 N44689 N44690 10
D44690 N44690 0 diode
R44691 N44690 N44691 10
D44691 N44691 0 diode
R44692 N44691 N44692 10
D44692 N44692 0 diode
R44693 N44692 N44693 10
D44693 N44693 0 diode
R44694 N44693 N44694 10
D44694 N44694 0 diode
R44695 N44694 N44695 10
D44695 N44695 0 diode
R44696 N44695 N44696 10
D44696 N44696 0 diode
R44697 N44696 N44697 10
D44697 N44697 0 diode
R44698 N44697 N44698 10
D44698 N44698 0 diode
R44699 N44698 N44699 10
D44699 N44699 0 diode
R44700 N44699 N44700 10
D44700 N44700 0 diode
R44701 N44700 N44701 10
D44701 N44701 0 diode
R44702 N44701 N44702 10
D44702 N44702 0 diode
R44703 N44702 N44703 10
D44703 N44703 0 diode
R44704 N44703 N44704 10
D44704 N44704 0 diode
R44705 N44704 N44705 10
D44705 N44705 0 diode
R44706 N44705 N44706 10
D44706 N44706 0 diode
R44707 N44706 N44707 10
D44707 N44707 0 diode
R44708 N44707 N44708 10
D44708 N44708 0 diode
R44709 N44708 N44709 10
D44709 N44709 0 diode
R44710 N44709 N44710 10
D44710 N44710 0 diode
R44711 N44710 N44711 10
D44711 N44711 0 diode
R44712 N44711 N44712 10
D44712 N44712 0 diode
R44713 N44712 N44713 10
D44713 N44713 0 diode
R44714 N44713 N44714 10
D44714 N44714 0 diode
R44715 N44714 N44715 10
D44715 N44715 0 diode
R44716 N44715 N44716 10
D44716 N44716 0 diode
R44717 N44716 N44717 10
D44717 N44717 0 diode
R44718 N44717 N44718 10
D44718 N44718 0 diode
R44719 N44718 N44719 10
D44719 N44719 0 diode
R44720 N44719 N44720 10
D44720 N44720 0 diode
R44721 N44720 N44721 10
D44721 N44721 0 diode
R44722 N44721 N44722 10
D44722 N44722 0 diode
R44723 N44722 N44723 10
D44723 N44723 0 diode
R44724 N44723 N44724 10
D44724 N44724 0 diode
R44725 N44724 N44725 10
D44725 N44725 0 diode
R44726 N44725 N44726 10
D44726 N44726 0 diode
R44727 N44726 N44727 10
D44727 N44727 0 diode
R44728 N44727 N44728 10
D44728 N44728 0 diode
R44729 N44728 N44729 10
D44729 N44729 0 diode
R44730 N44729 N44730 10
D44730 N44730 0 diode
R44731 N44730 N44731 10
D44731 N44731 0 diode
R44732 N44731 N44732 10
D44732 N44732 0 diode
R44733 N44732 N44733 10
D44733 N44733 0 diode
R44734 N44733 N44734 10
D44734 N44734 0 diode
R44735 N44734 N44735 10
D44735 N44735 0 diode
R44736 N44735 N44736 10
D44736 N44736 0 diode
R44737 N44736 N44737 10
D44737 N44737 0 diode
R44738 N44737 N44738 10
D44738 N44738 0 diode
R44739 N44738 N44739 10
D44739 N44739 0 diode
R44740 N44739 N44740 10
D44740 N44740 0 diode
R44741 N44740 N44741 10
D44741 N44741 0 diode
R44742 N44741 N44742 10
D44742 N44742 0 diode
R44743 N44742 N44743 10
D44743 N44743 0 diode
R44744 N44743 N44744 10
D44744 N44744 0 diode
R44745 N44744 N44745 10
D44745 N44745 0 diode
R44746 N44745 N44746 10
D44746 N44746 0 diode
R44747 N44746 N44747 10
D44747 N44747 0 diode
R44748 N44747 N44748 10
D44748 N44748 0 diode
R44749 N44748 N44749 10
D44749 N44749 0 diode
R44750 N44749 N44750 10
D44750 N44750 0 diode
R44751 N44750 N44751 10
D44751 N44751 0 diode
R44752 N44751 N44752 10
D44752 N44752 0 diode
R44753 N44752 N44753 10
D44753 N44753 0 diode
R44754 N44753 N44754 10
D44754 N44754 0 diode
R44755 N44754 N44755 10
D44755 N44755 0 diode
R44756 N44755 N44756 10
D44756 N44756 0 diode
R44757 N44756 N44757 10
D44757 N44757 0 diode
R44758 N44757 N44758 10
D44758 N44758 0 diode
R44759 N44758 N44759 10
D44759 N44759 0 diode
R44760 N44759 N44760 10
D44760 N44760 0 diode
R44761 N44760 N44761 10
D44761 N44761 0 diode
R44762 N44761 N44762 10
D44762 N44762 0 diode
R44763 N44762 N44763 10
D44763 N44763 0 diode
R44764 N44763 N44764 10
D44764 N44764 0 diode
R44765 N44764 N44765 10
D44765 N44765 0 diode
R44766 N44765 N44766 10
D44766 N44766 0 diode
R44767 N44766 N44767 10
D44767 N44767 0 diode
R44768 N44767 N44768 10
D44768 N44768 0 diode
R44769 N44768 N44769 10
D44769 N44769 0 diode
R44770 N44769 N44770 10
D44770 N44770 0 diode
R44771 N44770 N44771 10
D44771 N44771 0 diode
R44772 N44771 N44772 10
D44772 N44772 0 diode
R44773 N44772 N44773 10
D44773 N44773 0 diode
R44774 N44773 N44774 10
D44774 N44774 0 diode
R44775 N44774 N44775 10
D44775 N44775 0 diode
R44776 N44775 N44776 10
D44776 N44776 0 diode
R44777 N44776 N44777 10
D44777 N44777 0 diode
R44778 N44777 N44778 10
D44778 N44778 0 diode
R44779 N44778 N44779 10
D44779 N44779 0 diode
R44780 N44779 N44780 10
D44780 N44780 0 diode
R44781 N44780 N44781 10
D44781 N44781 0 diode
R44782 N44781 N44782 10
D44782 N44782 0 diode
R44783 N44782 N44783 10
D44783 N44783 0 diode
R44784 N44783 N44784 10
D44784 N44784 0 diode
R44785 N44784 N44785 10
D44785 N44785 0 diode
R44786 N44785 N44786 10
D44786 N44786 0 diode
R44787 N44786 N44787 10
D44787 N44787 0 diode
R44788 N44787 N44788 10
D44788 N44788 0 diode
R44789 N44788 N44789 10
D44789 N44789 0 diode
R44790 N44789 N44790 10
D44790 N44790 0 diode
R44791 N44790 N44791 10
D44791 N44791 0 diode
R44792 N44791 N44792 10
D44792 N44792 0 diode
R44793 N44792 N44793 10
D44793 N44793 0 diode
R44794 N44793 N44794 10
D44794 N44794 0 diode
R44795 N44794 N44795 10
D44795 N44795 0 diode
R44796 N44795 N44796 10
D44796 N44796 0 diode
R44797 N44796 N44797 10
D44797 N44797 0 diode
R44798 N44797 N44798 10
D44798 N44798 0 diode
R44799 N44798 N44799 10
D44799 N44799 0 diode
R44800 N44799 N44800 10
D44800 N44800 0 diode
R44801 N44800 N44801 10
D44801 N44801 0 diode
R44802 N44801 N44802 10
D44802 N44802 0 diode
R44803 N44802 N44803 10
D44803 N44803 0 diode
R44804 N44803 N44804 10
D44804 N44804 0 diode
R44805 N44804 N44805 10
D44805 N44805 0 diode
R44806 N44805 N44806 10
D44806 N44806 0 diode
R44807 N44806 N44807 10
D44807 N44807 0 diode
R44808 N44807 N44808 10
D44808 N44808 0 diode
R44809 N44808 N44809 10
D44809 N44809 0 diode
R44810 N44809 N44810 10
D44810 N44810 0 diode
R44811 N44810 N44811 10
D44811 N44811 0 diode
R44812 N44811 N44812 10
D44812 N44812 0 diode
R44813 N44812 N44813 10
D44813 N44813 0 diode
R44814 N44813 N44814 10
D44814 N44814 0 diode
R44815 N44814 N44815 10
D44815 N44815 0 diode
R44816 N44815 N44816 10
D44816 N44816 0 diode
R44817 N44816 N44817 10
D44817 N44817 0 diode
R44818 N44817 N44818 10
D44818 N44818 0 diode
R44819 N44818 N44819 10
D44819 N44819 0 diode
R44820 N44819 N44820 10
D44820 N44820 0 diode
R44821 N44820 N44821 10
D44821 N44821 0 diode
R44822 N44821 N44822 10
D44822 N44822 0 diode
R44823 N44822 N44823 10
D44823 N44823 0 diode
R44824 N44823 N44824 10
D44824 N44824 0 diode
R44825 N44824 N44825 10
D44825 N44825 0 diode
R44826 N44825 N44826 10
D44826 N44826 0 diode
R44827 N44826 N44827 10
D44827 N44827 0 diode
R44828 N44827 N44828 10
D44828 N44828 0 diode
R44829 N44828 N44829 10
D44829 N44829 0 diode
R44830 N44829 N44830 10
D44830 N44830 0 diode
R44831 N44830 N44831 10
D44831 N44831 0 diode
R44832 N44831 N44832 10
D44832 N44832 0 diode
R44833 N44832 N44833 10
D44833 N44833 0 diode
R44834 N44833 N44834 10
D44834 N44834 0 diode
R44835 N44834 N44835 10
D44835 N44835 0 diode
R44836 N44835 N44836 10
D44836 N44836 0 diode
R44837 N44836 N44837 10
D44837 N44837 0 diode
R44838 N44837 N44838 10
D44838 N44838 0 diode
R44839 N44838 N44839 10
D44839 N44839 0 diode
R44840 N44839 N44840 10
D44840 N44840 0 diode
R44841 N44840 N44841 10
D44841 N44841 0 diode
R44842 N44841 N44842 10
D44842 N44842 0 diode
R44843 N44842 N44843 10
D44843 N44843 0 diode
R44844 N44843 N44844 10
D44844 N44844 0 diode
R44845 N44844 N44845 10
D44845 N44845 0 diode
R44846 N44845 N44846 10
D44846 N44846 0 diode
R44847 N44846 N44847 10
D44847 N44847 0 diode
R44848 N44847 N44848 10
D44848 N44848 0 diode
R44849 N44848 N44849 10
D44849 N44849 0 diode
R44850 N44849 N44850 10
D44850 N44850 0 diode
R44851 N44850 N44851 10
D44851 N44851 0 diode
R44852 N44851 N44852 10
D44852 N44852 0 diode
R44853 N44852 N44853 10
D44853 N44853 0 diode
R44854 N44853 N44854 10
D44854 N44854 0 diode
R44855 N44854 N44855 10
D44855 N44855 0 diode
R44856 N44855 N44856 10
D44856 N44856 0 diode
R44857 N44856 N44857 10
D44857 N44857 0 diode
R44858 N44857 N44858 10
D44858 N44858 0 diode
R44859 N44858 N44859 10
D44859 N44859 0 diode
R44860 N44859 N44860 10
D44860 N44860 0 diode
R44861 N44860 N44861 10
D44861 N44861 0 diode
R44862 N44861 N44862 10
D44862 N44862 0 diode
R44863 N44862 N44863 10
D44863 N44863 0 diode
R44864 N44863 N44864 10
D44864 N44864 0 diode
R44865 N44864 N44865 10
D44865 N44865 0 diode
R44866 N44865 N44866 10
D44866 N44866 0 diode
R44867 N44866 N44867 10
D44867 N44867 0 diode
R44868 N44867 N44868 10
D44868 N44868 0 diode
R44869 N44868 N44869 10
D44869 N44869 0 diode
R44870 N44869 N44870 10
D44870 N44870 0 diode
R44871 N44870 N44871 10
D44871 N44871 0 diode
R44872 N44871 N44872 10
D44872 N44872 0 diode
R44873 N44872 N44873 10
D44873 N44873 0 diode
R44874 N44873 N44874 10
D44874 N44874 0 diode
R44875 N44874 N44875 10
D44875 N44875 0 diode
R44876 N44875 N44876 10
D44876 N44876 0 diode
R44877 N44876 N44877 10
D44877 N44877 0 diode
R44878 N44877 N44878 10
D44878 N44878 0 diode
R44879 N44878 N44879 10
D44879 N44879 0 diode
R44880 N44879 N44880 10
D44880 N44880 0 diode
R44881 N44880 N44881 10
D44881 N44881 0 diode
R44882 N44881 N44882 10
D44882 N44882 0 diode
R44883 N44882 N44883 10
D44883 N44883 0 diode
R44884 N44883 N44884 10
D44884 N44884 0 diode
R44885 N44884 N44885 10
D44885 N44885 0 diode
R44886 N44885 N44886 10
D44886 N44886 0 diode
R44887 N44886 N44887 10
D44887 N44887 0 diode
R44888 N44887 N44888 10
D44888 N44888 0 diode
R44889 N44888 N44889 10
D44889 N44889 0 diode
R44890 N44889 N44890 10
D44890 N44890 0 diode
R44891 N44890 N44891 10
D44891 N44891 0 diode
R44892 N44891 N44892 10
D44892 N44892 0 diode
R44893 N44892 N44893 10
D44893 N44893 0 diode
R44894 N44893 N44894 10
D44894 N44894 0 diode
R44895 N44894 N44895 10
D44895 N44895 0 diode
R44896 N44895 N44896 10
D44896 N44896 0 diode
R44897 N44896 N44897 10
D44897 N44897 0 diode
R44898 N44897 N44898 10
D44898 N44898 0 diode
R44899 N44898 N44899 10
D44899 N44899 0 diode
R44900 N44899 N44900 10
D44900 N44900 0 diode
R44901 N44900 N44901 10
D44901 N44901 0 diode
R44902 N44901 N44902 10
D44902 N44902 0 diode
R44903 N44902 N44903 10
D44903 N44903 0 diode
R44904 N44903 N44904 10
D44904 N44904 0 diode
R44905 N44904 N44905 10
D44905 N44905 0 diode
R44906 N44905 N44906 10
D44906 N44906 0 diode
R44907 N44906 N44907 10
D44907 N44907 0 diode
R44908 N44907 N44908 10
D44908 N44908 0 diode
R44909 N44908 N44909 10
D44909 N44909 0 diode
R44910 N44909 N44910 10
D44910 N44910 0 diode
R44911 N44910 N44911 10
D44911 N44911 0 diode
R44912 N44911 N44912 10
D44912 N44912 0 diode
R44913 N44912 N44913 10
D44913 N44913 0 diode
R44914 N44913 N44914 10
D44914 N44914 0 diode
R44915 N44914 N44915 10
D44915 N44915 0 diode
R44916 N44915 N44916 10
D44916 N44916 0 diode
R44917 N44916 N44917 10
D44917 N44917 0 diode
R44918 N44917 N44918 10
D44918 N44918 0 diode
R44919 N44918 N44919 10
D44919 N44919 0 diode
R44920 N44919 N44920 10
D44920 N44920 0 diode
R44921 N44920 N44921 10
D44921 N44921 0 diode
R44922 N44921 N44922 10
D44922 N44922 0 diode
R44923 N44922 N44923 10
D44923 N44923 0 diode
R44924 N44923 N44924 10
D44924 N44924 0 diode
R44925 N44924 N44925 10
D44925 N44925 0 diode
R44926 N44925 N44926 10
D44926 N44926 0 diode
R44927 N44926 N44927 10
D44927 N44927 0 diode
R44928 N44927 N44928 10
D44928 N44928 0 diode
R44929 N44928 N44929 10
D44929 N44929 0 diode
R44930 N44929 N44930 10
D44930 N44930 0 diode
R44931 N44930 N44931 10
D44931 N44931 0 diode
R44932 N44931 N44932 10
D44932 N44932 0 diode
R44933 N44932 N44933 10
D44933 N44933 0 diode
R44934 N44933 N44934 10
D44934 N44934 0 diode
R44935 N44934 N44935 10
D44935 N44935 0 diode
R44936 N44935 N44936 10
D44936 N44936 0 diode
R44937 N44936 N44937 10
D44937 N44937 0 diode
R44938 N44937 N44938 10
D44938 N44938 0 diode
R44939 N44938 N44939 10
D44939 N44939 0 diode
R44940 N44939 N44940 10
D44940 N44940 0 diode
R44941 N44940 N44941 10
D44941 N44941 0 diode
R44942 N44941 N44942 10
D44942 N44942 0 diode
R44943 N44942 N44943 10
D44943 N44943 0 diode
R44944 N44943 N44944 10
D44944 N44944 0 diode
R44945 N44944 N44945 10
D44945 N44945 0 diode
R44946 N44945 N44946 10
D44946 N44946 0 diode
R44947 N44946 N44947 10
D44947 N44947 0 diode
R44948 N44947 N44948 10
D44948 N44948 0 diode
R44949 N44948 N44949 10
D44949 N44949 0 diode
R44950 N44949 N44950 10
D44950 N44950 0 diode
R44951 N44950 N44951 10
D44951 N44951 0 diode
R44952 N44951 N44952 10
D44952 N44952 0 diode
R44953 N44952 N44953 10
D44953 N44953 0 diode
R44954 N44953 N44954 10
D44954 N44954 0 diode
R44955 N44954 N44955 10
D44955 N44955 0 diode
R44956 N44955 N44956 10
D44956 N44956 0 diode
R44957 N44956 N44957 10
D44957 N44957 0 diode
R44958 N44957 N44958 10
D44958 N44958 0 diode
R44959 N44958 N44959 10
D44959 N44959 0 diode
R44960 N44959 N44960 10
D44960 N44960 0 diode
R44961 N44960 N44961 10
D44961 N44961 0 diode
R44962 N44961 N44962 10
D44962 N44962 0 diode
R44963 N44962 N44963 10
D44963 N44963 0 diode
R44964 N44963 N44964 10
D44964 N44964 0 diode
R44965 N44964 N44965 10
D44965 N44965 0 diode
R44966 N44965 N44966 10
D44966 N44966 0 diode
R44967 N44966 N44967 10
D44967 N44967 0 diode
R44968 N44967 N44968 10
D44968 N44968 0 diode
R44969 N44968 N44969 10
D44969 N44969 0 diode
R44970 N44969 N44970 10
D44970 N44970 0 diode
R44971 N44970 N44971 10
D44971 N44971 0 diode
R44972 N44971 N44972 10
D44972 N44972 0 diode
R44973 N44972 N44973 10
D44973 N44973 0 diode
R44974 N44973 N44974 10
D44974 N44974 0 diode
R44975 N44974 N44975 10
D44975 N44975 0 diode
R44976 N44975 N44976 10
D44976 N44976 0 diode
R44977 N44976 N44977 10
D44977 N44977 0 diode
R44978 N44977 N44978 10
D44978 N44978 0 diode
R44979 N44978 N44979 10
D44979 N44979 0 diode
R44980 N44979 N44980 10
D44980 N44980 0 diode
R44981 N44980 N44981 10
D44981 N44981 0 diode
R44982 N44981 N44982 10
D44982 N44982 0 diode
R44983 N44982 N44983 10
D44983 N44983 0 diode
R44984 N44983 N44984 10
D44984 N44984 0 diode
R44985 N44984 N44985 10
D44985 N44985 0 diode
R44986 N44985 N44986 10
D44986 N44986 0 diode
R44987 N44986 N44987 10
D44987 N44987 0 diode
R44988 N44987 N44988 10
D44988 N44988 0 diode
R44989 N44988 N44989 10
D44989 N44989 0 diode
R44990 N44989 N44990 10
D44990 N44990 0 diode
R44991 N44990 N44991 10
D44991 N44991 0 diode
R44992 N44991 N44992 10
D44992 N44992 0 diode
R44993 N44992 N44993 10
D44993 N44993 0 diode
R44994 N44993 N44994 10
D44994 N44994 0 diode
R44995 N44994 N44995 10
D44995 N44995 0 diode
R44996 N44995 N44996 10
D44996 N44996 0 diode
R44997 N44996 N44997 10
D44997 N44997 0 diode
R44998 N44997 N44998 10
D44998 N44998 0 diode
R44999 N44998 N44999 10
D44999 N44999 0 diode
R45000 N44999 N45000 10
D45000 N45000 0 diode
R45001 N45000 N45001 10
D45001 N45001 0 diode
R45002 N45001 N45002 10
D45002 N45002 0 diode
R45003 N45002 N45003 10
D45003 N45003 0 diode
R45004 N45003 N45004 10
D45004 N45004 0 diode
R45005 N45004 N45005 10
D45005 N45005 0 diode
R45006 N45005 N45006 10
D45006 N45006 0 diode
R45007 N45006 N45007 10
D45007 N45007 0 diode
R45008 N45007 N45008 10
D45008 N45008 0 diode
R45009 N45008 N45009 10
D45009 N45009 0 diode
R45010 N45009 N45010 10
D45010 N45010 0 diode
R45011 N45010 N45011 10
D45011 N45011 0 diode
R45012 N45011 N45012 10
D45012 N45012 0 diode
R45013 N45012 N45013 10
D45013 N45013 0 diode
R45014 N45013 N45014 10
D45014 N45014 0 diode
R45015 N45014 N45015 10
D45015 N45015 0 diode
R45016 N45015 N45016 10
D45016 N45016 0 diode
R45017 N45016 N45017 10
D45017 N45017 0 diode
R45018 N45017 N45018 10
D45018 N45018 0 diode
R45019 N45018 N45019 10
D45019 N45019 0 diode
R45020 N45019 N45020 10
D45020 N45020 0 diode
R45021 N45020 N45021 10
D45021 N45021 0 diode
R45022 N45021 N45022 10
D45022 N45022 0 diode
R45023 N45022 N45023 10
D45023 N45023 0 diode
R45024 N45023 N45024 10
D45024 N45024 0 diode
R45025 N45024 N45025 10
D45025 N45025 0 diode
R45026 N45025 N45026 10
D45026 N45026 0 diode
R45027 N45026 N45027 10
D45027 N45027 0 diode
R45028 N45027 N45028 10
D45028 N45028 0 diode
R45029 N45028 N45029 10
D45029 N45029 0 diode
R45030 N45029 N45030 10
D45030 N45030 0 diode
R45031 N45030 N45031 10
D45031 N45031 0 diode
R45032 N45031 N45032 10
D45032 N45032 0 diode
R45033 N45032 N45033 10
D45033 N45033 0 diode
R45034 N45033 N45034 10
D45034 N45034 0 diode
R45035 N45034 N45035 10
D45035 N45035 0 diode
R45036 N45035 N45036 10
D45036 N45036 0 diode
R45037 N45036 N45037 10
D45037 N45037 0 diode
R45038 N45037 N45038 10
D45038 N45038 0 diode
R45039 N45038 N45039 10
D45039 N45039 0 diode
R45040 N45039 N45040 10
D45040 N45040 0 diode
R45041 N45040 N45041 10
D45041 N45041 0 diode
R45042 N45041 N45042 10
D45042 N45042 0 diode
R45043 N45042 N45043 10
D45043 N45043 0 diode
R45044 N45043 N45044 10
D45044 N45044 0 diode
R45045 N45044 N45045 10
D45045 N45045 0 diode
R45046 N45045 N45046 10
D45046 N45046 0 diode
R45047 N45046 N45047 10
D45047 N45047 0 diode
R45048 N45047 N45048 10
D45048 N45048 0 diode
R45049 N45048 N45049 10
D45049 N45049 0 diode
R45050 N45049 N45050 10
D45050 N45050 0 diode
R45051 N45050 N45051 10
D45051 N45051 0 diode
R45052 N45051 N45052 10
D45052 N45052 0 diode
R45053 N45052 N45053 10
D45053 N45053 0 diode
R45054 N45053 N45054 10
D45054 N45054 0 diode
R45055 N45054 N45055 10
D45055 N45055 0 diode
R45056 N45055 N45056 10
D45056 N45056 0 diode
R45057 N45056 N45057 10
D45057 N45057 0 diode
R45058 N45057 N45058 10
D45058 N45058 0 diode
R45059 N45058 N45059 10
D45059 N45059 0 diode
R45060 N45059 N45060 10
D45060 N45060 0 diode
R45061 N45060 N45061 10
D45061 N45061 0 diode
R45062 N45061 N45062 10
D45062 N45062 0 diode
R45063 N45062 N45063 10
D45063 N45063 0 diode
R45064 N45063 N45064 10
D45064 N45064 0 diode
R45065 N45064 N45065 10
D45065 N45065 0 diode
R45066 N45065 N45066 10
D45066 N45066 0 diode
R45067 N45066 N45067 10
D45067 N45067 0 diode
R45068 N45067 N45068 10
D45068 N45068 0 diode
R45069 N45068 N45069 10
D45069 N45069 0 diode
R45070 N45069 N45070 10
D45070 N45070 0 diode
R45071 N45070 N45071 10
D45071 N45071 0 diode
R45072 N45071 N45072 10
D45072 N45072 0 diode
R45073 N45072 N45073 10
D45073 N45073 0 diode
R45074 N45073 N45074 10
D45074 N45074 0 diode
R45075 N45074 N45075 10
D45075 N45075 0 diode
R45076 N45075 N45076 10
D45076 N45076 0 diode
R45077 N45076 N45077 10
D45077 N45077 0 diode
R45078 N45077 N45078 10
D45078 N45078 0 diode
R45079 N45078 N45079 10
D45079 N45079 0 diode
R45080 N45079 N45080 10
D45080 N45080 0 diode
R45081 N45080 N45081 10
D45081 N45081 0 diode
R45082 N45081 N45082 10
D45082 N45082 0 diode
R45083 N45082 N45083 10
D45083 N45083 0 diode
R45084 N45083 N45084 10
D45084 N45084 0 diode
R45085 N45084 N45085 10
D45085 N45085 0 diode
R45086 N45085 N45086 10
D45086 N45086 0 diode
R45087 N45086 N45087 10
D45087 N45087 0 diode
R45088 N45087 N45088 10
D45088 N45088 0 diode
R45089 N45088 N45089 10
D45089 N45089 0 diode
R45090 N45089 N45090 10
D45090 N45090 0 diode
R45091 N45090 N45091 10
D45091 N45091 0 diode
R45092 N45091 N45092 10
D45092 N45092 0 diode
R45093 N45092 N45093 10
D45093 N45093 0 diode
R45094 N45093 N45094 10
D45094 N45094 0 diode
R45095 N45094 N45095 10
D45095 N45095 0 diode
R45096 N45095 N45096 10
D45096 N45096 0 diode
R45097 N45096 N45097 10
D45097 N45097 0 diode
R45098 N45097 N45098 10
D45098 N45098 0 diode
R45099 N45098 N45099 10
D45099 N45099 0 diode
R45100 N45099 N45100 10
D45100 N45100 0 diode
R45101 N45100 N45101 10
D45101 N45101 0 diode
R45102 N45101 N45102 10
D45102 N45102 0 diode
R45103 N45102 N45103 10
D45103 N45103 0 diode
R45104 N45103 N45104 10
D45104 N45104 0 diode
R45105 N45104 N45105 10
D45105 N45105 0 diode
R45106 N45105 N45106 10
D45106 N45106 0 diode
R45107 N45106 N45107 10
D45107 N45107 0 diode
R45108 N45107 N45108 10
D45108 N45108 0 diode
R45109 N45108 N45109 10
D45109 N45109 0 diode
R45110 N45109 N45110 10
D45110 N45110 0 diode
R45111 N45110 N45111 10
D45111 N45111 0 diode
R45112 N45111 N45112 10
D45112 N45112 0 diode
R45113 N45112 N45113 10
D45113 N45113 0 diode
R45114 N45113 N45114 10
D45114 N45114 0 diode
R45115 N45114 N45115 10
D45115 N45115 0 diode
R45116 N45115 N45116 10
D45116 N45116 0 diode
R45117 N45116 N45117 10
D45117 N45117 0 diode
R45118 N45117 N45118 10
D45118 N45118 0 diode
R45119 N45118 N45119 10
D45119 N45119 0 diode
R45120 N45119 N45120 10
D45120 N45120 0 diode
R45121 N45120 N45121 10
D45121 N45121 0 diode
R45122 N45121 N45122 10
D45122 N45122 0 diode
R45123 N45122 N45123 10
D45123 N45123 0 diode
R45124 N45123 N45124 10
D45124 N45124 0 diode
R45125 N45124 N45125 10
D45125 N45125 0 diode
R45126 N45125 N45126 10
D45126 N45126 0 diode
R45127 N45126 N45127 10
D45127 N45127 0 diode
R45128 N45127 N45128 10
D45128 N45128 0 diode
R45129 N45128 N45129 10
D45129 N45129 0 diode
R45130 N45129 N45130 10
D45130 N45130 0 diode
R45131 N45130 N45131 10
D45131 N45131 0 diode
R45132 N45131 N45132 10
D45132 N45132 0 diode
R45133 N45132 N45133 10
D45133 N45133 0 diode
R45134 N45133 N45134 10
D45134 N45134 0 diode
R45135 N45134 N45135 10
D45135 N45135 0 diode
R45136 N45135 N45136 10
D45136 N45136 0 diode
R45137 N45136 N45137 10
D45137 N45137 0 diode
R45138 N45137 N45138 10
D45138 N45138 0 diode
R45139 N45138 N45139 10
D45139 N45139 0 diode
R45140 N45139 N45140 10
D45140 N45140 0 diode
R45141 N45140 N45141 10
D45141 N45141 0 diode
R45142 N45141 N45142 10
D45142 N45142 0 diode
R45143 N45142 N45143 10
D45143 N45143 0 diode
R45144 N45143 N45144 10
D45144 N45144 0 diode
R45145 N45144 N45145 10
D45145 N45145 0 diode
R45146 N45145 N45146 10
D45146 N45146 0 diode
R45147 N45146 N45147 10
D45147 N45147 0 diode
R45148 N45147 N45148 10
D45148 N45148 0 diode
R45149 N45148 N45149 10
D45149 N45149 0 diode
R45150 N45149 N45150 10
D45150 N45150 0 diode
R45151 N45150 N45151 10
D45151 N45151 0 diode
R45152 N45151 N45152 10
D45152 N45152 0 diode
R45153 N45152 N45153 10
D45153 N45153 0 diode
R45154 N45153 N45154 10
D45154 N45154 0 diode
R45155 N45154 N45155 10
D45155 N45155 0 diode
R45156 N45155 N45156 10
D45156 N45156 0 diode
R45157 N45156 N45157 10
D45157 N45157 0 diode
R45158 N45157 N45158 10
D45158 N45158 0 diode
R45159 N45158 N45159 10
D45159 N45159 0 diode
R45160 N45159 N45160 10
D45160 N45160 0 diode
R45161 N45160 N45161 10
D45161 N45161 0 diode
R45162 N45161 N45162 10
D45162 N45162 0 diode
R45163 N45162 N45163 10
D45163 N45163 0 diode
R45164 N45163 N45164 10
D45164 N45164 0 diode
R45165 N45164 N45165 10
D45165 N45165 0 diode
R45166 N45165 N45166 10
D45166 N45166 0 diode
R45167 N45166 N45167 10
D45167 N45167 0 diode
R45168 N45167 N45168 10
D45168 N45168 0 diode
R45169 N45168 N45169 10
D45169 N45169 0 diode
R45170 N45169 N45170 10
D45170 N45170 0 diode
R45171 N45170 N45171 10
D45171 N45171 0 diode
R45172 N45171 N45172 10
D45172 N45172 0 diode
R45173 N45172 N45173 10
D45173 N45173 0 diode
R45174 N45173 N45174 10
D45174 N45174 0 diode
R45175 N45174 N45175 10
D45175 N45175 0 diode
R45176 N45175 N45176 10
D45176 N45176 0 diode
R45177 N45176 N45177 10
D45177 N45177 0 diode
R45178 N45177 N45178 10
D45178 N45178 0 diode
R45179 N45178 N45179 10
D45179 N45179 0 diode
R45180 N45179 N45180 10
D45180 N45180 0 diode
R45181 N45180 N45181 10
D45181 N45181 0 diode
R45182 N45181 N45182 10
D45182 N45182 0 diode
R45183 N45182 N45183 10
D45183 N45183 0 diode
R45184 N45183 N45184 10
D45184 N45184 0 diode
R45185 N45184 N45185 10
D45185 N45185 0 diode
R45186 N45185 N45186 10
D45186 N45186 0 diode
R45187 N45186 N45187 10
D45187 N45187 0 diode
R45188 N45187 N45188 10
D45188 N45188 0 diode
R45189 N45188 N45189 10
D45189 N45189 0 diode
R45190 N45189 N45190 10
D45190 N45190 0 diode
R45191 N45190 N45191 10
D45191 N45191 0 diode
R45192 N45191 N45192 10
D45192 N45192 0 diode
R45193 N45192 N45193 10
D45193 N45193 0 diode
R45194 N45193 N45194 10
D45194 N45194 0 diode
R45195 N45194 N45195 10
D45195 N45195 0 diode
R45196 N45195 N45196 10
D45196 N45196 0 diode
R45197 N45196 N45197 10
D45197 N45197 0 diode
R45198 N45197 N45198 10
D45198 N45198 0 diode
R45199 N45198 N45199 10
D45199 N45199 0 diode
R45200 N45199 N45200 10
D45200 N45200 0 diode
R45201 N45200 N45201 10
D45201 N45201 0 diode
R45202 N45201 N45202 10
D45202 N45202 0 diode
R45203 N45202 N45203 10
D45203 N45203 0 diode
R45204 N45203 N45204 10
D45204 N45204 0 diode
R45205 N45204 N45205 10
D45205 N45205 0 diode
R45206 N45205 N45206 10
D45206 N45206 0 diode
R45207 N45206 N45207 10
D45207 N45207 0 diode
R45208 N45207 N45208 10
D45208 N45208 0 diode
R45209 N45208 N45209 10
D45209 N45209 0 diode
R45210 N45209 N45210 10
D45210 N45210 0 diode
R45211 N45210 N45211 10
D45211 N45211 0 diode
R45212 N45211 N45212 10
D45212 N45212 0 diode
R45213 N45212 N45213 10
D45213 N45213 0 diode
R45214 N45213 N45214 10
D45214 N45214 0 diode
R45215 N45214 N45215 10
D45215 N45215 0 diode
R45216 N45215 N45216 10
D45216 N45216 0 diode
R45217 N45216 N45217 10
D45217 N45217 0 diode
R45218 N45217 N45218 10
D45218 N45218 0 diode
R45219 N45218 N45219 10
D45219 N45219 0 diode
R45220 N45219 N45220 10
D45220 N45220 0 diode
R45221 N45220 N45221 10
D45221 N45221 0 diode
R45222 N45221 N45222 10
D45222 N45222 0 diode
R45223 N45222 N45223 10
D45223 N45223 0 diode
R45224 N45223 N45224 10
D45224 N45224 0 diode
R45225 N45224 N45225 10
D45225 N45225 0 diode
R45226 N45225 N45226 10
D45226 N45226 0 diode
R45227 N45226 N45227 10
D45227 N45227 0 diode
R45228 N45227 N45228 10
D45228 N45228 0 diode
R45229 N45228 N45229 10
D45229 N45229 0 diode
R45230 N45229 N45230 10
D45230 N45230 0 diode
R45231 N45230 N45231 10
D45231 N45231 0 diode
R45232 N45231 N45232 10
D45232 N45232 0 diode
R45233 N45232 N45233 10
D45233 N45233 0 diode
R45234 N45233 N45234 10
D45234 N45234 0 diode
R45235 N45234 N45235 10
D45235 N45235 0 diode
R45236 N45235 N45236 10
D45236 N45236 0 diode
R45237 N45236 N45237 10
D45237 N45237 0 diode
R45238 N45237 N45238 10
D45238 N45238 0 diode
R45239 N45238 N45239 10
D45239 N45239 0 diode
R45240 N45239 N45240 10
D45240 N45240 0 diode
R45241 N45240 N45241 10
D45241 N45241 0 diode
R45242 N45241 N45242 10
D45242 N45242 0 diode
R45243 N45242 N45243 10
D45243 N45243 0 diode
R45244 N45243 N45244 10
D45244 N45244 0 diode
R45245 N45244 N45245 10
D45245 N45245 0 diode
R45246 N45245 N45246 10
D45246 N45246 0 diode
R45247 N45246 N45247 10
D45247 N45247 0 diode
R45248 N45247 N45248 10
D45248 N45248 0 diode
R45249 N45248 N45249 10
D45249 N45249 0 diode
R45250 N45249 N45250 10
D45250 N45250 0 diode
R45251 N45250 N45251 10
D45251 N45251 0 diode
R45252 N45251 N45252 10
D45252 N45252 0 diode
R45253 N45252 N45253 10
D45253 N45253 0 diode
R45254 N45253 N45254 10
D45254 N45254 0 diode
R45255 N45254 N45255 10
D45255 N45255 0 diode
R45256 N45255 N45256 10
D45256 N45256 0 diode
R45257 N45256 N45257 10
D45257 N45257 0 diode
R45258 N45257 N45258 10
D45258 N45258 0 diode
R45259 N45258 N45259 10
D45259 N45259 0 diode
R45260 N45259 N45260 10
D45260 N45260 0 diode
R45261 N45260 N45261 10
D45261 N45261 0 diode
R45262 N45261 N45262 10
D45262 N45262 0 diode
R45263 N45262 N45263 10
D45263 N45263 0 diode
R45264 N45263 N45264 10
D45264 N45264 0 diode
R45265 N45264 N45265 10
D45265 N45265 0 diode
R45266 N45265 N45266 10
D45266 N45266 0 diode
R45267 N45266 N45267 10
D45267 N45267 0 diode
R45268 N45267 N45268 10
D45268 N45268 0 diode
R45269 N45268 N45269 10
D45269 N45269 0 diode
R45270 N45269 N45270 10
D45270 N45270 0 diode
R45271 N45270 N45271 10
D45271 N45271 0 diode
R45272 N45271 N45272 10
D45272 N45272 0 diode
R45273 N45272 N45273 10
D45273 N45273 0 diode
R45274 N45273 N45274 10
D45274 N45274 0 diode
R45275 N45274 N45275 10
D45275 N45275 0 diode
R45276 N45275 N45276 10
D45276 N45276 0 diode
R45277 N45276 N45277 10
D45277 N45277 0 diode
R45278 N45277 N45278 10
D45278 N45278 0 diode
R45279 N45278 N45279 10
D45279 N45279 0 diode
R45280 N45279 N45280 10
D45280 N45280 0 diode
R45281 N45280 N45281 10
D45281 N45281 0 diode
R45282 N45281 N45282 10
D45282 N45282 0 diode
R45283 N45282 N45283 10
D45283 N45283 0 diode
R45284 N45283 N45284 10
D45284 N45284 0 diode
R45285 N45284 N45285 10
D45285 N45285 0 diode
R45286 N45285 N45286 10
D45286 N45286 0 diode
R45287 N45286 N45287 10
D45287 N45287 0 diode
R45288 N45287 N45288 10
D45288 N45288 0 diode
R45289 N45288 N45289 10
D45289 N45289 0 diode
R45290 N45289 N45290 10
D45290 N45290 0 diode
R45291 N45290 N45291 10
D45291 N45291 0 diode
R45292 N45291 N45292 10
D45292 N45292 0 diode
R45293 N45292 N45293 10
D45293 N45293 0 diode
R45294 N45293 N45294 10
D45294 N45294 0 diode
R45295 N45294 N45295 10
D45295 N45295 0 diode
R45296 N45295 N45296 10
D45296 N45296 0 diode
R45297 N45296 N45297 10
D45297 N45297 0 diode
R45298 N45297 N45298 10
D45298 N45298 0 diode
R45299 N45298 N45299 10
D45299 N45299 0 diode
R45300 N45299 N45300 10
D45300 N45300 0 diode
R45301 N45300 N45301 10
D45301 N45301 0 diode
R45302 N45301 N45302 10
D45302 N45302 0 diode
R45303 N45302 N45303 10
D45303 N45303 0 diode
R45304 N45303 N45304 10
D45304 N45304 0 diode
R45305 N45304 N45305 10
D45305 N45305 0 diode
R45306 N45305 N45306 10
D45306 N45306 0 diode
R45307 N45306 N45307 10
D45307 N45307 0 diode
R45308 N45307 N45308 10
D45308 N45308 0 diode
R45309 N45308 N45309 10
D45309 N45309 0 diode
R45310 N45309 N45310 10
D45310 N45310 0 diode
R45311 N45310 N45311 10
D45311 N45311 0 diode
R45312 N45311 N45312 10
D45312 N45312 0 diode
R45313 N45312 N45313 10
D45313 N45313 0 diode
R45314 N45313 N45314 10
D45314 N45314 0 diode
R45315 N45314 N45315 10
D45315 N45315 0 diode
R45316 N45315 N45316 10
D45316 N45316 0 diode
R45317 N45316 N45317 10
D45317 N45317 0 diode
R45318 N45317 N45318 10
D45318 N45318 0 diode
R45319 N45318 N45319 10
D45319 N45319 0 diode
R45320 N45319 N45320 10
D45320 N45320 0 diode
R45321 N45320 N45321 10
D45321 N45321 0 diode
R45322 N45321 N45322 10
D45322 N45322 0 diode
R45323 N45322 N45323 10
D45323 N45323 0 diode
R45324 N45323 N45324 10
D45324 N45324 0 diode
R45325 N45324 N45325 10
D45325 N45325 0 diode
R45326 N45325 N45326 10
D45326 N45326 0 diode
R45327 N45326 N45327 10
D45327 N45327 0 diode
R45328 N45327 N45328 10
D45328 N45328 0 diode
R45329 N45328 N45329 10
D45329 N45329 0 diode
R45330 N45329 N45330 10
D45330 N45330 0 diode
R45331 N45330 N45331 10
D45331 N45331 0 diode
R45332 N45331 N45332 10
D45332 N45332 0 diode
R45333 N45332 N45333 10
D45333 N45333 0 diode
R45334 N45333 N45334 10
D45334 N45334 0 diode
R45335 N45334 N45335 10
D45335 N45335 0 diode
R45336 N45335 N45336 10
D45336 N45336 0 diode
R45337 N45336 N45337 10
D45337 N45337 0 diode
R45338 N45337 N45338 10
D45338 N45338 0 diode
R45339 N45338 N45339 10
D45339 N45339 0 diode
R45340 N45339 N45340 10
D45340 N45340 0 diode
R45341 N45340 N45341 10
D45341 N45341 0 diode
R45342 N45341 N45342 10
D45342 N45342 0 diode
R45343 N45342 N45343 10
D45343 N45343 0 diode
R45344 N45343 N45344 10
D45344 N45344 0 diode
R45345 N45344 N45345 10
D45345 N45345 0 diode
R45346 N45345 N45346 10
D45346 N45346 0 diode
R45347 N45346 N45347 10
D45347 N45347 0 diode
R45348 N45347 N45348 10
D45348 N45348 0 diode
R45349 N45348 N45349 10
D45349 N45349 0 diode
R45350 N45349 N45350 10
D45350 N45350 0 diode
R45351 N45350 N45351 10
D45351 N45351 0 diode
R45352 N45351 N45352 10
D45352 N45352 0 diode
R45353 N45352 N45353 10
D45353 N45353 0 diode
R45354 N45353 N45354 10
D45354 N45354 0 diode
R45355 N45354 N45355 10
D45355 N45355 0 diode
R45356 N45355 N45356 10
D45356 N45356 0 diode
R45357 N45356 N45357 10
D45357 N45357 0 diode
R45358 N45357 N45358 10
D45358 N45358 0 diode
R45359 N45358 N45359 10
D45359 N45359 0 diode
R45360 N45359 N45360 10
D45360 N45360 0 diode
R45361 N45360 N45361 10
D45361 N45361 0 diode
R45362 N45361 N45362 10
D45362 N45362 0 diode
R45363 N45362 N45363 10
D45363 N45363 0 diode
R45364 N45363 N45364 10
D45364 N45364 0 diode
R45365 N45364 N45365 10
D45365 N45365 0 diode
R45366 N45365 N45366 10
D45366 N45366 0 diode
R45367 N45366 N45367 10
D45367 N45367 0 diode
R45368 N45367 N45368 10
D45368 N45368 0 diode
R45369 N45368 N45369 10
D45369 N45369 0 diode
R45370 N45369 N45370 10
D45370 N45370 0 diode
R45371 N45370 N45371 10
D45371 N45371 0 diode
R45372 N45371 N45372 10
D45372 N45372 0 diode
R45373 N45372 N45373 10
D45373 N45373 0 diode
R45374 N45373 N45374 10
D45374 N45374 0 diode
R45375 N45374 N45375 10
D45375 N45375 0 diode
R45376 N45375 N45376 10
D45376 N45376 0 diode
R45377 N45376 N45377 10
D45377 N45377 0 diode
R45378 N45377 N45378 10
D45378 N45378 0 diode
R45379 N45378 N45379 10
D45379 N45379 0 diode
R45380 N45379 N45380 10
D45380 N45380 0 diode
R45381 N45380 N45381 10
D45381 N45381 0 diode
R45382 N45381 N45382 10
D45382 N45382 0 diode
R45383 N45382 N45383 10
D45383 N45383 0 diode
R45384 N45383 N45384 10
D45384 N45384 0 diode
R45385 N45384 N45385 10
D45385 N45385 0 diode
R45386 N45385 N45386 10
D45386 N45386 0 diode
R45387 N45386 N45387 10
D45387 N45387 0 diode
R45388 N45387 N45388 10
D45388 N45388 0 diode
R45389 N45388 N45389 10
D45389 N45389 0 diode
R45390 N45389 N45390 10
D45390 N45390 0 diode
R45391 N45390 N45391 10
D45391 N45391 0 diode
R45392 N45391 N45392 10
D45392 N45392 0 diode
R45393 N45392 N45393 10
D45393 N45393 0 diode
R45394 N45393 N45394 10
D45394 N45394 0 diode
R45395 N45394 N45395 10
D45395 N45395 0 diode
R45396 N45395 N45396 10
D45396 N45396 0 diode
R45397 N45396 N45397 10
D45397 N45397 0 diode
R45398 N45397 N45398 10
D45398 N45398 0 diode
R45399 N45398 N45399 10
D45399 N45399 0 diode
R45400 N45399 N45400 10
D45400 N45400 0 diode
R45401 N45400 N45401 10
D45401 N45401 0 diode
R45402 N45401 N45402 10
D45402 N45402 0 diode
R45403 N45402 N45403 10
D45403 N45403 0 diode
R45404 N45403 N45404 10
D45404 N45404 0 diode
R45405 N45404 N45405 10
D45405 N45405 0 diode
R45406 N45405 N45406 10
D45406 N45406 0 diode
R45407 N45406 N45407 10
D45407 N45407 0 diode
R45408 N45407 N45408 10
D45408 N45408 0 diode
R45409 N45408 N45409 10
D45409 N45409 0 diode
R45410 N45409 N45410 10
D45410 N45410 0 diode
R45411 N45410 N45411 10
D45411 N45411 0 diode
R45412 N45411 N45412 10
D45412 N45412 0 diode
R45413 N45412 N45413 10
D45413 N45413 0 diode
R45414 N45413 N45414 10
D45414 N45414 0 diode
R45415 N45414 N45415 10
D45415 N45415 0 diode
R45416 N45415 N45416 10
D45416 N45416 0 diode
R45417 N45416 N45417 10
D45417 N45417 0 diode
R45418 N45417 N45418 10
D45418 N45418 0 diode
R45419 N45418 N45419 10
D45419 N45419 0 diode
R45420 N45419 N45420 10
D45420 N45420 0 diode
R45421 N45420 N45421 10
D45421 N45421 0 diode
R45422 N45421 N45422 10
D45422 N45422 0 diode
R45423 N45422 N45423 10
D45423 N45423 0 diode
R45424 N45423 N45424 10
D45424 N45424 0 diode
R45425 N45424 N45425 10
D45425 N45425 0 diode
R45426 N45425 N45426 10
D45426 N45426 0 diode
R45427 N45426 N45427 10
D45427 N45427 0 diode
R45428 N45427 N45428 10
D45428 N45428 0 diode
R45429 N45428 N45429 10
D45429 N45429 0 diode
R45430 N45429 N45430 10
D45430 N45430 0 diode
R45431 N45430 N45431 10
D45431 N45431 0 diode
R45432 N45431 N45432 10
D45432 N45432 0 diode
R45433 N45432 N45433 10
D45433 N45433 0 diode
R45434 N45433 N45434 10
D45434 N45434 0 diode
R45435 N45434 N45435 10
D45435 N45435 0 diode
R45436 N45435 N45436 10
D45436 N45436 0 diode
R45437 N45436 N45437 10
D45437 N45437 0 diode
R45438 N45437 N45438 10
D45438 N45438 0 diode
R45439 N45438 N45439 10
D45439 N45439 0 diode
R45440 N45439 N45440 10
D45440 N45440 0 diode
R45441 N45440 N45441 10
D45441 N45441 0 diode
R45442 N45441 N45442 10
D45442 N45442 0 diode
R45443 N45442 N45443 10
D45443 N45443 0 diode
R45444 N45443 N45444 10
D45444 N45444 0 diode
R45445 N45444 N45445 10
D45445 N45445 0 diode
R45446 N45445 N45446 10
D45446 N45446 0 diode
R45447 N45446 N45447 10
D45447 N45447 0 diode
R45448 N45447 N45448 10
D45448 N45448 0 diode
R45449 N45448 N45449 10
D45449 N45449 0 diode
R45450 N45449 N45450 10
D45450 N45450 0 diode
R45451 N45450 N45451 10
D45451 N45451 0 diode
R45452 N45451 N45452 10
D45452 N45452 0 diode
R45453 N45452 N45453 10
D45453 N45453 0 diode
R45454 N45453 N45454 10
D45454 N45454 0 diode
R45455 N45454 N45455 10
D45455 N45455 0 diode
R45456 N45455 N45456 10
D45456 N45456 0 diode
R45457 N45456 N45457 10
D45457 N45457 0 diode
R45458 N45457 N45458 10
D45458 N45458 0 diode
R45459 N45458 N45459 10
D45459 N45459 0 diode
R45460 N45459 N45460 10
D45460 N45460 0 diode
R45461 N45460 N45461 10
D45461 N45461 0 diode
R45462 N45461 N45462 10
D45462 N45462 0 diode
R45463 N45462 N45463 10
D45463 N45463 0 diode
R45464 N45463 N45464 10
D45464 N45464 0 diode
R45465 N45464 N45465 10
D45465 N45465 0 diode
R45466 N45465 N45466 10
D45466 N45466 0 diode
R45467 N45466 N45467 10
D45467 N45467 0 diode
R45468 N45467 N45468 10
D45468 N45468 0 diode
R45469 N45468 N45469 10
D45469 N45469 0 diode
R45470 N45469 N45470 10
D45470 N45470 0 diode
R45471 N45470 N45471 10
D45471 N45471 0 diode
R45472 N45471 N45472 10
D45472 N45472 0 diode
R45473 N45472 N45473 10
D45473 N45473 0 diode
R45474 N45473 N45474 10
D45474 N45474 0 diode
R45475 N45474 N45475 10
D45475 N45475 0 diode
R45476 N45475 N45476 10
D45476 N45476 0 diode
R45477 N45476 N45477 10
D45477 N45477 0 diode
R45478 N45477 N45478 10
D45478 N45478 0 diode
R45479 N45478 N45479 10
D45479 N45479 0 diode
R45480 N45479 N45480 10
D45480 N45480 0 diode
R45481 N45480 N45481 10
D45481 N45481 0 diode
R45482 N45481 N45482 10
D45482 N45482 0 diode
R45483 N45482 N45483 10
D45483 N45483 0 diode
R45484 N45483 N45484 10
D45484 N45484 0 diode
R45485 N45484 N45485 10
D45485 N45485 0 diode
R45486 N45485 N45486 10
D45486 N45486 0 diode
R45487 N45486 N45487 10
D45487 N45487 0 diode
R45488 N45487 N45488 10
D45488 N45488 0 diode
R45489 N45488 N45489 10
D45489 N45489 0 diode
R45490 N45489 N45490 10
D45490 N45490 0 diode
R45491 N45490 N45491 10
D45491 N45491 0 diode
R45492 N45491 N45492 10
D45492 N45492 0 diode
R45493 N45492 N45493 10
D45493 N45493 0 diode
R45494 N45493 N45494 10
D45494 N45494 0 diode
R45495 N45494 N45495 10
D45495 N45495 0 diode
R45496 N45495 N45496 10
D45496 N45496 0 diode
R45497 N45496 N45497 10
D45497 N45497 0 diode
R45498 N45497 N45498 10
D45498 N45498 0 diode
R45499 N45498 N45499 10
D45499 N45499 0 diode
R45500 N45499 N45500 10
D45500 N45500 0 diode
R45501 N45500 N45501 10
D45501 N45501 0 diode
R45502 N45501 N45502 10
D45502 N45502 0 diode
R45503 N45502 N45503 10
D45503 N45503 0 diode
R45504 N45503 N45504 10
D45504 N45504 0 diode
R45505 N45504 N45505 10
D45505 N45505 0 diode
R45506 N45505 N45506 10
D45506 N45506 0 diode
R45507 N45506 N45507 10
D45507 N45507 0 diode
R45508 N45507 N45508 10
D45508 N45508 0 diode
R45509 N45508 N45509 10
D45509 N45509 0 diode
R45510 N45509 N45510 10
D45510 N45510 0 diode
R45511 N45510 N45511 10
D45511 N45511 0 diode
R45512 N45511 N45512 10
D45512 N45512 0 diode
R45513 N45512 N45513 10
D45513 N45513 0 diode
R45514 N45513 N45514 10
D45514 N45514 0 diode
R45515 N45514 N45515 10
D45515 N45515 0 diode
R45516 N45515 N45516 10
D45516 N45516 0 diode
R45517 N45516 N45517 10
D45517 N45517 0 diode
R45518 N45517 N45518 10
D45518 N45518 0 diode
R45519 N45518 N45519 10
D45519 N45519 0 diode
R45520 N45519 N45520 10
D45520 N45520 0 diode
R45521 N45520 N45521 10
D45521 N45521 0 diode
R45522 N45521 N45522 10
D45522 N45522 0 diode
R45523 N45522 N45523 10
D45523 N45523 0 diode
R45524 N45523 N45524 10
D45524 N45524 0 diode
R45525 N45524 N45525 10
D45525 N45525 0 diode
R45526 N45525 N45526 10
D45526 N45526 0 diode
R45527 N45526 N45527 10
D45527 N45527 0 diode
R45528 N45527 N45528 10
D45528 N45528 0 diode
R45529 N45528 N45529 10
D45529 N45529 0 diode
R45530 N45529 N45530 10
D45530 N45530 0 diode
R45531 N45530 N45531 10
D45531 N45531 0 diode
R45532 N45531 N45532 10
D45532 N45532 0 diode
R45533 N45532 N45533 10
D45533 N45533 0 diode
R45534 N45533 N45534 10
D45534 N45534 0 diode
R45535 N45534 N45535 10
D45535 N45535 0 diode
R45536 N45535 N45536 10
D45536 N45536 0 diode
R45537 N45536 N45537 10
D45537 N45537 0 diode
R45538 N45537 N45538 10
D45538 N45538 0 diode
R45539 N45538 N45539 10
D45539 N45539 0 diode
R45540 N45539 N45540 10
D45540 N45540 0 diode
R45541 N45540 N45541 10
D45541 N45541 0 diode
R45542 N45541 N45542 10
D45542 N45542 0 diode
R45543 N45542 N45543 10
D45543 N45543 0 diode
R45544 N45543 N45544 10
D45544 N45544 0 diode
R45545 N45544 N45545 10
D45545 N45545 0 diode
R45546 N45545 N45546 10
D45546 N45546 0 diode
R45547 N45546 N45547 10
D45547 N45547 0 diode
R45548 N45547 N45548 10
D45548 N45548 0 diode
R45549 N45548 N45549 10
D45549 N45549 0 diode
R45550 N45549 N45550 10
D45550 N45550 0 diode
R45551 N45550 N45551 10
D45551 N45551 0 diode
R45552 N45551 N45552 10
D45552 N45552 0 diode
R45553 N45552 N45553 10
D45553 N45553 0 diode
R45554 N45553 N45554 10
D45554 N45554 0 diode
R45555 N45554 N45555 10
D45555 N45555 0 diode
R45556 N45555 N45556 10
D45556 N45556 0 diode
R45557 N45556 N45557 10
D45557 N45557 0 diode
R45558 N45557 N45558 10
D45558 N45558 0 diode
R45559 N45558 N45559 10
D45559 N45559 0 diode
R45560 N45559 N45560 10
D45560 N45560 0 diode
R45561 N45560 N45561 10
D45561 N45561 0 diode
R45562 N45561 N45562 10
D45562 N45562 0 diode
R45563 N45562 N45563 10
D45563 N45563 0 diode
R45564 N45563 N45564 10
D45564 N45564 0 diode
R45565 N45564 N45565 10
D45565 N45565 0 diode
R45566 N45565 N45566 10
D45566 N45566 0 diode
R45567 N45566 N45567 10
D45567 N45567 0 diode
R45568 N45567 N45568 10
D45568 N45568 0 diode
R45569 N45568 N45569 10
D45569 N45569 0 diode
R45570 N45569 N45570 10
D45570 N45570 0 diode
R45571 N45570 N45571 10
D45571 N45571 0 diode
R45572 N45571 N45572 10
D45572 N45572 0 diode
R45573 N45572 N45573 10
D45573 N45573 0 diode
R45574 N45573 N45574 10
D45574 N45574 0 diode
R45575 N45574 N45575 10
D45575 N45575 0 diode
R45576 N45575 N45576 10
D45576 N45576 0 diode
R45577 N45576 N45577 10
D45577 N45577 0 diode
R45578 N45577 N45578 10
D45578 N45578 0 diode
R45579 N45578 N45579 10
D45579 N45579 0 diode
R45580 N45579 N45580 10
D45580 N45580 0 diode
R45581 N45580 N45581 10
D45581 N45581 0 diode
R45582 N45581 N45582 10
D45582 N45582 0 diode
R45583 N45582 N45583 10
D45583 N45583 0 diode
R45584 N45583 N45584 10
D45584 N45584 0 diode
R45585 N45584 N45585 10
D45585 N45585 0 diode
R45586 N45585 N45586 10
D45586 N45586 0 diode
R45587 N45586 N45587 10
D45587 N45587 0 diode
R45588 N45587 N45588 10
D45588 N45588 0 diode
R45589 N45588 N45589 10
D45589 N45589 0 diode
R45590 N45589 N45590 10
D45590 N45590 0 diode
R45591 N45590 N45591 10
D45591 N45591 0 diode
R45592 N45591 N45592 10
D45592 N45592 0 diode
R45593 N45592 N45593 10
D45593 N45593 0 diode
R45594 N45593 N45594 10
D45594 N45594 0 diode
R45595 N45594 N45595 10
D45595 N45595 0 diode
R45596 N45595 N45596 10
D45596 N45596 0 diode
R45597 N45596 N45597 10
D45597 N45597 0 diode
R45598 N45597 N45598 10
D45598 N45598 0 diode
R45599 N45598 N45599 10
D45599 N45599 0 diode
R45600 N45599 N45600 10
D45600 N45600 0 diode
R45601 N45600 N45601 10
D45601 N45601 0 diode
R45602 N45601 N45602 10
D45602 N45602 0 diode
R45603 N45602 N45603 10
D45603 N45603 0 diode
R45604 N45603 N45604 10
D45604 N45604 0 diode
R45605 N45604 N45605 10
D45605 N45605 0 diode
R45606 N45605 N45606 10
D45606 N45606 0 diode
R45607 N45606 N45607 10
D45607 N45607 0 diode
R45608 N45607 N45608 10
D45608 N45608 0 diode
R45609 N45608 N45609 10
D45609 N45609 0 diode
R45610 N45609 N45610 10
D45610 N45610 0 diode
R45611 N45610 N45611 10
D45611 N45611 0 diode
R45612 N45611 N45612 10
D45612 N45612 0 diode
R45613 N45612 N45613 10
D45613 N45613 0 diode
R45614 N45613 N45614 10
D45614 N45614 0 diode
R45615 N45614 N45615 10
D45615 N45615 0 diode
R45616 N45615 N45616 10
D45616 N45616 0 diode
R45617 N45616 N45617 10
D45617 N45617 0 diode
R45618 N45617 N45618 10
D45618 N45618 0 diode
R45619 N45618 N45619 10
D45619 N45619 0 diode
R45620 N45619 N45620 10
D45620 N45620 0 diode
R45621 N45620 N45621 10
D45621 N45621 0 diode
R45622 N45621 N45622 10
D45622 N45622 0 diode
R45623 N45622 N45623 10
D45623 N45623 0 diode
R45624 N45623 N45624 10
D45624 N45624 0 diode
R45625 N45624 N45625 10
D45625 N45625 0 diode
R45626 N45625 N45626 10
D45626 N45626 0 diode
R45627 N45626 N45627 10
D45627 N45627 0 diode
R45628 N45627 N45628 10
D45628 N45628 0 diode
R45629 N45628 N45629 10
D45629 N45629 0 diode
R45630 N45629 N45630 10
D45630 N45630 0 diode
R45631 N45630 N45631 10
D45631 N45631 0 diode
R45632 N45631 N45632 10
D45632 N45632 0 diode
R45633 N45632 N45633 10
D45633 N45633 0 diode
R45634 N45633 N45634 10
D45634 N45634 0 diode
R45635 N45634 N45635 10
D45635 N45635 0 diode
R45636 N45635 N45636 10
D45636 N45636 0 diode
R45637 N45636 N45637 10
D45637 N45637 0 diode
R45638 N45637 N45638 10
D45638 N45638 0 diode
R45639 N45638 N45639 10
D45639 N45639 0 diode
R45640 N45639 N45640 10
D45640 N45640 0 diode
R45641 N45640 N45641 10
D45641 N45641 0 diode
R45642 N45641 N45642 10
D45642 N45642 0 diode
R45643 N45642 N45643 10
D45643 N45643 0 diode
R45644 N45643 N45644 10
D45644 N45644 0 diode
R45645 N45644 N45645 10
D45645 N45645 0 diode
R45646 N45645 N45646 10
D45646 N45646 0 diode
R45647 N45646 N45647 10
D45647 N45647 0 diode
R45648 N45647 N45648 10
D45648 N45648 0 diode
R45649 N45648 N45649 10
D45649 N45649 0 diode
R45650 N45649 N45650 10
D45650 N45650 0 diode
R45651 N45650 N45651 10
D45651 N45651 0 diode
R45652 N45651 N45652 10
D45652 N45652 0 diode
R45653 N45652 N45653 10
D45653 N45653 0 diode
R45654 N45653 N45654 10
D45654 N45654 0 diode
R45655 N45654 N45655 10
D45655 N45655 0 diode
R45656 N45655 N45656 10
D45656 N45656 0 diode
R45657 N45656 N45657 10
D45657 N45657 0 diode
R45658 N45657 N45658 10
D45658 N45658 0 diode
R45659 N45658 N45659 10
D45659 N45659 0 diode
R45660 N45659 N45660 10
D45660 N45660 0 diode
R45661 N45660 N45661 10
D45661 N45661 0 diode
R45662 N45661 N45662 10
D45662 N45662 0 diode
R45663 N45662 N45663 10
D45663 N45663 0 diode
R45664 N45663 N45664 10
D45664 N45664 0 diode
R45665 N45664 N45665 10
D45665 N45665 0 diode
R45666 N45665 N45666 10
D45666 N45666 0 diode
R45667 N45666 N45667 10
D45667 N45667 0 diode
R45668 N45667 N45668 10
D45668 N45668 0 diode
R45669 N45668 N45669 10
D45669 N45669 0 diode
R45670 N45669 N45670 10
D45670 N45670 0 diode
R45671 N45670 N45671 10
D45671 N45671 0 diode
R45672 N45671 N45672 10
D45672 N45672 0 diode
R45673 N45672 N45673 10
D45673 N45673 0 diode
R45674 N45673 N45674 10
D45674 N45674 0 diode
R45675 N45674 N45675 10
D45675 N45675 0 diode
R45676 N45675 N45676 10
D45676 N45676 0 diode
R45677 N45676 N45677 10
D45677 N45677 0 diode
R45678 N45677 N45678 10
D45678 N45678 0 diode
R45679 N45678 N45679 10
D45679 N45679 0 diode
R45680 N45679 N45680 10
D45680 N45680 0 diode
R45681 N45680 N45681 10
D45681 N45681 0 diode
R45682 N45681 N45682 10
D45682 N45682 0 diode
R45683 N45682 N45683 10
D45683 N45683 0 diode
R45684 N45683 N45684 10
D45684 N45684 0 diode
R45685 N45684 N45685 10
D45685 N45685 0 diode
R45686 N45685 N45686 10
D45686 N45686 0 diode
R45687 N45686 N45687 10
D45687 N45687 0 diode
R45688 N45687 N45688 10
D45688 N45688 0 diode
R45689 N45688 N45689 10
D45689 N45689 0 diode
R45690 N45689 N45690 10
D45690 N45690 0 diode
R45691 N45690 N45691 10
D45691 N45691 0 diode
R45692 N45691 N45692 10
D45692 N45692 0 diode
R45693 N45692 N45693 10
D45693 N45693 0 diode
R45694 N45693 N45694 10
D45694 N45694 0 diode
R45695 N45694 N45695 10
D45695 N45695 0 diode
R45696 N45695 N45696 10
D45696 N45696 0 diode
R45697 N45696 N45697 10
D45697 N45697 0 diode
R45698 N45697 N45698 10
D45698 N45698 0 diode
R45699 N45698 N45699 10
D45699 N45699 0 diode
R45700 N45699 N45700 10
D45700 N45700 0 diode
R45701 N45700 N45701 10
D45701 N45701 0 diode
R45702 N45701 N45702 10
D45702 N45702 0 diode
R45703 N45702 N45703 10
D45703 N45703 0 diode
R45704 N45703 N45704 10
D45704 N45704 0 diode
R45705 N45704 N45705 10
D45705 N45705 0 diode
R45706 N45705 N45706 10
D45706 N45706 0 diode
R45707 N45706 N45707 10
D45707 N45707 0 diode
R45708 N45707 N45708 10
D45708 N45708 0 diode
R45709 N45708 N45709 10
D45709 N45709 0 diode
R45710 N45709 N45710 10
D45710 N45710 0 diode
R45711 N45710 N45711 10
D45711 N45711 0 diode
R45712 N45711 N45712 10
D45712 N45712 0 diode
R45713 N45712 N45713 10
D45713 N45713 0 diode
R45714 N45713 N45714 10
D45714 N45714 0 diode
R45715 N45714 N45715 10
D45715 N45715 0 diode
R45716 N45715 N45716 10
D45716 N45716 0 diode
R45717 N45716 N45717 10
D45717 N45717 0 diode
R45718 N45717 N45718 10
D45718 N45718 0 diode
R45719 N45718 N45719 10
D45719 N45719 0 diode
R45720 N45719 N45720 10
D45720 N45720 0 diode
R45721 N45720 N45721 10
D45721 N45721 0 diode
R45722 N45721 N45722 10
D45722 N45722 0 diode
R45723 N45722 N45723 10
D45723 N45723 0 diode
R45724 N45723 N45724 10
D45724 N45724 0 diode
R45725 N45724 N45725 10
D45725 N45725 0 diode
R45726 N45725 N45726 10
D45726 N45726 0 diode
R45727 N45726 N45727 10
D45727 N45727 0 diode
R45728 N45727 N45728 10
D45728 N45728 0 diode
R45729 N45728 N45729 10
D45729 N45729 0 diode
R45730 N45729 N45730 10
D45730 N45730 0 diode
R45731 N45730 N45731 10
D45731 N45731 0 diode
R45732 N45731 N45732 10
D45732 N45732 0 diode
R45733 N45732 N45733 10
D45733 N45733 0 diode
R45734 N45733 N45734 10
D45734 N45734 0 diode
R45735 N45734 N45735 10
D45735 N45735 0 diode
R45736 N45735 N45736 10
D45736 N45736 0 diode
R45737 N45736 N45737 10
D45737 N45737 0 diode
R45738 N45737 N45738 10
D45738 N45738 0 diode
R45739 N45738 N45739 10
D45739 N45739 0 diode
R45740 N45739 N45740 10
D45740 N45740 0 diode
R45741 N45740 N45741 10
D45741 N45741 0 diode
R45742 N45741 N45742 10
D45742 N45742 0 diode
R45743 N45742 N45743 10
D45743 N45743 0 diode
R45744 N45743 N45744 10
D45744 N45744 0 diode
R45745 N45744 N45745 10
D45745 N45745 0 diode
R45746 N45745 N45746 10
D45746 N45746 0 diode
R45747 N45746 N45747 10
D45747 N45747 0 diode
R45748 N45747 N45748 10
D45748 N45748 0 diode
R45749 N45748 N45749 10
D45749 N45749 0 diode
R45750 N45749 N45750 10
D45750 N45750 0 diode
R45751 N45750 N45751 10
D45751 N45751 0 diode
R45752 N45751 N45752 10
D45752 N45752 0 diode
R45753 N45752 N45753 10
D45753 N45753 0 diode
R45754 N45753 N45754 10
D45754 N45754 0 diode
R45755 N45754 N45755 10
D45755 N45755 0 diode
R45756 N45755 N45756 10
D45756 N45756 0 diode
R45757 N45756 N45757 10
D45757 N45757 0 diode
R45758 N45757 N45758 10
D45758 N45758 0 diode
R45759 N45758 N45759 10
D45759 N45759 0 diode
R45760 N45759 N45760 10
D45760 N45760 0 diode
R45761 N45760 N45761 10
D45761 N45761 0 diode
R45762 N45761 N45762 10
D45762 N45762 0 diode
R45763 N45762 N45763 10
D45763 N45763 0 diode
R45764 N45763 N45764 10
D45764 N45764 0 diode
R45765 N45764 N45765 10
D45765 N45765 0 diode
R45766 N45765 N45766 10
D45766 N45766 0 diode
R45767 N45766 N45767 10
D45767 N45767 0 diode
R45768 N45767 N45768 10
D45768 N45768 0 diode
R45769 N45768 N45769 10
D45769 N45769 0 diode
R45770 N45769 N45770 10
D45770 N45770 0 diode
R45771 N45770 N45771 10
D45771 N45771 0 diode
R45772 N45771 N45772 10
D45772 N45772 0 diode
R45773 N45772 N45773 10
D45773 N45773 0 diode
R45774 N45773 N45774 10
D45774 N45774 0 diode
R45775 N45774 N45775 10
D45775 N45775 0 diode
R45776 N45775 N45776 10
D45776 N45776 0 diode
R45777 N45776 N45777 10
D45777 N45777 0 diode
R45778 N45777 N45778 10
D45778 N45778 0 diode
R45779 N45778 N45779 10
D45779 N45779 0 diode
R45780 N45779 N45780 10
D45780 N45780 0 diode
R45781 N45780 N45781 10
D45781 N45781 0 diode
R45782 N45781 N45782 10
D45782 N45782 0 diode
R45783 N45782 N45783 10
D45783 N45783 0 diode
R45784 N45783 N45784 10
D45784 N45784 0 diode
R45785 N45784 N45785 10
D45785 N45785 0 diode
R45786 N45785 N45786 10
D45786 N45786 0 diode
R45787 N45786 N45787 10
D45787 N45787 0 diode
R45788 N45787 N45788 10
D45788 N45788 0 diode
R45789 N45788 N45789 10
D45789 N45789 0 diode
R45790 N45789 N45790 10
D45790 N45790 0 diode
R45791 N45790 N45791 10
D45791 N45791 0 diode
R45792 N45791 N45792 10
D45792 N45792 0 diode
R45793 N45792 N45793 10
D45793 N45793 0 diode
R45794 N45793 N45794 10
D45794 N45794 0 diode
R45795 N45794 N45795 10
D45795 N45795 0 diode
R45796 N45795 N45796 10
D45796 N45796 0 diode
R45797 N45796 N45797 10
D45797 N45797 0 diode
R45798 N45797 N45798 10
D45798 N45798 0 diode
R45799 N45798 N45799 10
D45799 N45799 0 diode
R45800 N45799 N45800 10
D45800 N45800 0 diode
R45801 N45800 N45801 10
D45801 N45801 0 diode
R45802 N45801 N45802 10
D45802 N45802 0 diode
R45803 N45802 N45803 10
D45803 N45803 0 diode
R45804 N45803 N45804 10
D45804 N45804 0 diode
R45805 N45804 N45805 10
D45805 N45805 0 diode
R45806 N45805 N45806 10
D45806 N45806 0 diode
R45807 N45806 N45807 10
D45807 N45807 0 diode
R45808 N45807 N45808 10
D45808 N45808 0 diode
R45809 N45808 N45809 10
D45809 N45809 0 diode
R45810 N45809 N45810 10
D45810 N45810 0 diode
R45811 N45810 N45811 10
D45811 N45811 0 diode
R45812 N45811 N45812 10
D45812 N45812 0 diode
R45813 N45812 N45813 10
D45813 N45813 0 diode
R45814 N45813 N45814 10
D45814 N45814 0 diode
R45815 N45814 N45815 10
D45815 N45815 0 diode
R45816 N45815 N45816 10
D45816 N45816 0 diode
R45817 N45816 N45817 10
D45817 N45817 0 diode
R45818 N45817 N45818 10
D45818 N45818 0 diode
R45819 N45818 N45819 10
D45819 N45819 0 diode
R45820 N45819 N45820 10
D45820 N45820 0 diode
R45821 N45820 N45821 10
D45821 N45821 0 diode
R45822 N45821 N45822 10
D45822 N45822 0 diode
R45823 N45822 N45823 10
D45823 N45823 0 diode
R45824 N45823 N45824 10
D45824 N45824 0 diode
R45825 N45824 N45825 10
D45825 N45825 0 diode
R45826 N45825 N45826 10
D45826 N45826 0 diode
R45827 N45826 N45827 10
D45827 N45827 0 diode
R45828 N45827 N45828 10
D45828 N45828 0 diode
R45829 N45828 N45829 10
D45829 N45829 0 diode
R45830 N45829 N45830 10
D45830 N45830 0 diode
R45831 N45830 N45831 10
D45831 N45831 0 diode
R45832 N45831 N45832 10
D45832 N45832 0 diode
R45833 N45832 N45833 10
D45833 N45833 0 diode
R45834 N45833 N45834 10
D45834 N45834 0 diode
R45835 N45834 N45835 10
D45835 N45835 0 diode
R45836 N45835 N45836 10
D45836 N45836 0 diode
R45837 N45836 N45837 10
D45837 N45837 0 diode
R45838 N45837 N45838 10
D45838 N45838 0 diode
R45839 N45838 N45839 10
D45839 N45839 0 diode
R45840 N45839 N45840 10
D45840 N45840 0 diode
R45841 N45840 N45841 10
D45841 N45841 0 diode
R45842 N45841 N45842 10
D45842 N45842 0 diode
R45843 N45842 N45843 10
D45843 N45843 0 diode
R45844 N45843 N45844 10
D45844 N45844 0 diode
R45845 N45844 N45845 10
D45845 N45845 0 diode
R45846 N45845 N45846 10
D45846 N45846 0 diode
R45847 N45846 N45847 10
D45847 N45847 0 diode
R45848 N45847 N45848 10
D45848 N45848 0 diode
R45849 N45848 N45849 10
D45849 N45849 0 diode
R45850 N45849 N45850 10
D45850 N45850 0 diode
R45851 N45850 N45851 10
D45851 N45851 0 diode
R45852 N45851 N45852 10
D45852 N45852 0 diode
R45853 N45852 N45853 10
D45853 N45853 0 diode
R45854 N45853 N45854 10
D45854 N45854 0 diode
R45855 N45854 N45855 10
D45855 N45855 0 diode
R45856 N45855 N45856 10
D45856 N45856 0 diode
R45857 N45856 N45857 10
D45857 N45857 0 diode
R45858 N45857 N45858 10
D45858 N45858 0 diode
R45859 N45858 N45859 10
D45859 N45859 0 diode
R45860 N45859 N45860 10
D45860 N45860 0 diode
R45861 N45860 N45861 10
D45861 N45861 0 diode
R45862 N45861 N45862 10
D45862 N45862 0 diode
R45863 N45862 N45863 10
D45863 N45863 0 diode
R45864 N45863 N45864 10
D45864 N45864 0 diode
R45865 N45864 N45865 10
D45865 N45865 0 diode
R45866 N45865 N45866 10
D45866 N45866 0 diode
R45867 N45866 N45867 10
D45867 N45867 0 diode
R45868 N45867 N45868 10
D45868 N45868 0 diode
R45869 N45868 N45869 10
D45869 N45869 0 diode
R45870 N45869 N45870 10
D45870 N45870 0 diode
R45871 N45870 N45871 10
D45871 N45871 0 diode
R45872 N45871 N45872 10
D45872 N45872 0 diode
R45873 N45872 N45873 10
D45873 N45873 0 diode
R45874 N45873 N45874 10
D45874 N45874 0 diode
R45875 N45874 N45875 10
D45875 N45875 0 diode
R45876 N45875 N45876 10
D45876 N45876 0 diode
R45877 N45876 N45877 10
D45877 N45877 0 diode
R45878 N45877 N45878 10
D45878 N45878 0 diode
R45879 N45878 N45879 10
D45879 N45879 0 diode
R45880 N45879 N45880 10
D45880 N45880 0 diode
R45881 N45880 N45881 10
D45881 N45881 0 diode
R45882 N45881 N45882 10
D45882 N45882 0 diode
R45883 N45882 N45883 10
D45883 N45883 0 diode
R45884 N45883 N45884 10
D45884 N45884 0 diode
R45885 N45884 N45885 10
D45885 N45885 0 diode
R45886 N45885 N45886 10
D45886 N45886 0 diode
R45887 N45886 N45887 10
D45887 N45887 0 diode
R45888 N45887 N45888 10
D45888 N45888 0 diode
R45889 N45888 N45889 10
D45889 N45889 0 diode
R45890 N45889 N45890 10
D45890 N45890 0 diode
R45891 N45890 N45891 10
D45891 N45891 0 diode
R45892 N45891 N45892 10
D45892 N45892 0 diode
R45893 N45892 N45893 10
D45893 N45893 0 diode
R45894 N45893 N45894 10
D45894 N45894 0 diode
R45895 N45894 N45895 10
D45895 N45895 0 diode
R45896 N45895 N45896 10
D45896 N45896 0 diode
R45897 N45896 N45897 10
D45897 N45897 0 diode
R45898 N45897 N45898 10
D45898 N45898 0 diode
R45899 N45898 N45899 10
D45899 N45899 0 diode
R45900 N45899 N45900 10
D45900 N45900 0 diode
R45901 N45900 N45901 10
D45901 N45901 0 diode
R45902 N45901 N45902 10
D45902 N45902 0 diode
R45903 N45902 N45903 10
D45903 N45903 0 diode
R45904 N45903 N45904 10
D45904 N45904 0 diode
R45905 N45904 N45905 10
D45905 N45905 0 diode
R45906 N45905 N45906 10
D45906 N45906 0 diode
R45907 N45906 N45907 10
D45907 N45907 0 diode
R45908 N45907 N45908 10
D45908 N45908 0 diode
R45909 N45908 N45909 10
D45909 N45909 0 diode
R45910 N45909 N45910 10
D45910 N45910 0 diode
R45911 N45910 N45911 10
D45911 N45911 0 diode
R45912 N45911 N45912 10
D45912 N45912 0 diode
R45913 N45912 N45913 10
D45913 N45913 0 diode
R45914 N45913 N45914 10
D45914 N45914 0 diode
R45915 N45914 N45915 10
D45915 N45915 0 diode
R45916 N45915 N45916 10
D45916 N45916 0 diode
R45917 N45916 N45917 10
D45917 N45917 0 diode
R45918 N45917 N45918 10
D45918 N45918 0 diode
R45919 N45918 N45919 10
D45919 N45919 0 diode
R45920 N45919 N45920 10
D45920 N45920 0 diode
R45921 N45920 N45921 10
D45921 N45921 0 diode
R45922 N45921 N45922 10
D45922 N45922 0 diode
R45923 N45922 N45923 10
D45923 N45923 0 diode
R45924 N45923 N45924 10
D45924 N45924 0 diode
R45925 N45924 N45925 10
D45925 N45925 0 diode
R45926 N45925 N45926 10
D45926 N45926 0 diode
R45927 N45926 N45927 10
D45927 N45927 0 diode
R45928 N45927 N45928 10
D45928 N45928 0 diode
R45929 N45928 N45929 10
D45929 N45929 0 diode
R45930 N45929 N45930 10
D45930 N45930 0 diode
R45931 N45930 N45931 10
D45931 N45931 0 diode
R45932 N45931 N45932 10
D45932 N45932 0 diode
R45933 N45932 N45933 10
D45933 N45933 0 diode
R45934 N45933 N45934 10
D45934 N45934 0 diode
R45935 N45934 N45935 10
D45935 N45935 0 diode
R45936 N45935 N45936 10
D45936 N45936 0 diode
R45937 N45936 N45937 10
D45937 N45937 0 diode
R45938 N45937 N45938 10
D45938 N45938 0 diode
R45939 N45938 N45939 10
D45939 N45939 0 diode
R45940 N45939 N45940 10
D45940 N45940 0 diode
R45941 N45940 N45941 10
D45941 N45941 0 diode
R45942 N45941 N45942 10
D45942 N45942 0 diode
R45943 N45942 N45943 10
D45943 N45943 0 diode
R45944 N45943 N45944 10
D45944 N45944 0 diode
R45945 N45944 N45945 10
D45945 N45945 0 diode
R45946 N45945 N45946 10
D45946 N45946 0 diode
R45947 N45946 N45947 10
D45947 N45947 0 diode
R45948 N45947 N45948 10
D45948 N45948 0 diode
R45949 N45948 N45949 10
D45949 N45949 0 diode
R45950 N45949 N45950 10
D45950 N45950 0 diode
R45951 N45950 N45951 10
D45951 N45951 0 diode
R45952 N45951 N45952 10
D45952 N45952 0 diode
R45953 N45952 N45953 10
D45953 N45953 0 diode
R45954 N45953 N45954 10
D45954 N45954 0 diode
R45955 N45954 N45955 10
D45955 N45955 0 diode
R45956 N45955 N45956 10
D45956 N45956 0 diode
R45957 N45956 N45957 10
D45957 N45957 0 diode
R45958 N45957 N45958 10
D45958 N45958 0 diode
R45959 N45958 N45959 10
D45959 N45959 0 diode
R45960 N45959 N45960 10
D45960 N45960 0 diode
R45961 N45960 N45961 10
D45961 N45961 0 diode
R45962 N45961 N45962 10
D45962 N45962 0 diode
R45963 N45962 N45963 10
D45963 N45963 0 diode
R45964 N45963 N45964 10
D45964 N45964 0 diode
R45965 N45964 N45965 10
D45965 N45965 0 diode
R45966 N45965 N45966 10
D45966 N45966 0 diode
R45967 N45966 N45967 10
D45967 N45967 0 diode
R45968 N45967 N45968 10
D45968 N45968 0 diode
R45969 N45968 N45969 10
D45969 N45969 0 diode
R45970 N45969 N45970 10
D45970 N45970 0 diode
R45971 N45970 N45971 10
D45971 N45971 0 diode
R45972 N45971 N45972 10
D45972 N45972 0 diode
R45973 N45972 N45973 10
D45973 N45973 0 diode
R45974 N45973 N45974 10
D45974 N45974 0 diode
R45975 N45974 N45975 10
D45975 N45975 0 diode
R45976 N45975 N45976 10
D45976 N45976 0 diode
R45977 N45976 N45977 10
D45977 N45977 0 diode
R45978 N45977 N45978 10
D45978 N45978 0 diode
R45979 N45978 N45979 10
D45979 N45979 0 diode
R45980 N45979 N45980 10
D45980 N45980 0 diode
R45981 N45980 N45981 10
D45981 N45981 0 diode
R45982 N45981 N45982 10
D45982 N45982 0 diode
R45983 N45982 N45983 10
D45983 N45983 0 diode
R45984 N45983 N45984 10
D45984 N45984 0 diode
R45985 N45984 N45985 10
D45985 N45985 0 diode
R45986 N45985 N45986 10
D45986 N45986 0 diode
R45987 N45986 N45987 10
D45987 N45987 0 diode
R45988 N45987 N45988 10
D45988 N45988 0 diode
R45989 N45988 N45989 10
D45989 N45989 0 diode
R45990 N45989 N45990 10
D45990 N45990 0 diode
R45991 N45990 N45991 10
D45991 N45991 0 diode
R45992 N45991 N45992 10
D45992 N45992 0 diode
R45993 N45992 N45993 10
D45993 N45993 0 diode
R45994 N45993 N45994 10
D45994 N45994 0 diode
R45995 N45994 N45995 10
D45995 N45995 0 diode
R45996 N45995 N45996 10
D45996 N45996 0 diode
R45997 N45996 N45997 10
D45997 N45997 0 diode
R45998 N45997 N45998 10
D45998 N45998 0 diode
R45999 N45998 N45999 10
D45999 N45999 0 diode
R46000 N45999 N46000 10
D46000 N46000 0 diode
R46001 N46000 N46001 10
D46001 N46001 0 diode
R46002 N46001 N46002 10
D46002 N46002 0 diode
R46003 N46002 N46003 10
D46003 N46003 0 diode
R46004 N46003 N46004 10
D46004 N46004 0 diode
R46005 N46004 N46005 10
D46005 N46005 0 diode
R46006 N46005 N46006 10
D46006 N46006 0 diode
R46007 N46006 N46007 10
D46007 N46007 0 diode
R46008 N46007 N46008 10
D46008 N46008 0 diode
R46009 N46008 N46009 10
D46009 N46009 0 diode
R46010 N46009 N46010 10
D46010 N46010 0 diode
R46011 N46010 N46011 10
D46011 N46011 0 diode
R46012 N46011 N46012 10
D46012 N46012 0 diode
R46013 N46012 N46013 10
D46013 N46013 0 diode
R46014 N46013 N46014 10
D46014 N46014 0 diode
R46015 N46014 N46015 10
D46015 N46015 0 diode
R46016 N46015 N46016 10
D46016 N46016 0 diode
R46017 N46016 N46017 10
D46017 N46017 0 diode
R46018 N46017 N46018 10
D46018 N46018 0 diode
R46019 N46018 N46019 10
D46019 N46019 0 diode
R46020 N46019 N46020 10
D46020 N46020 0 diode
R46021 N46020 N46021 10
D46021 N46021 0 diode
R46022 N46021 N46022 10
D46022 N46022 0 diode
R46023 N46022 N46023 10
D46023 N46023 0 diode
R46024 N46023 N46024 10
D46024 N46024 0 diode
R46025 N46024 N46025 10
D46025 N46025 0 diode
R46026 N46025 N46026 10
D46026 N46026 0 diode
R46027 N46026 N46027 10
D46027 N46027 0 diode
R46028 N46027 N46028 10
D46028 N46028 0 diode
R46029 N46028 N46029 10
D46029 N46029 0 diode
R46030 N46029 N46030 10
D46030 N46030 0 diode
R46031 N46030 N46031 10
D46031 N46031 0 diode
R46032 N46031 N46032 10
D46032 N46032 0 diode
R46033 N46032 N46033 10
D46033 N46033 0 diode
R46034 N46033 N46034 10
D46034 N46034 0 diode
R46035 N46034 N46035 10
D46035 N46035 0 diode
R46036 N46035 N46036 10
D46036 N46036 0 diode
R46037 N46036 N46037 10
D46037 N46037 0 diode
R46038 N46037 N46038 10
D46038 N46038 0 diode
R46039 N46038 N46039 10
D46039 N46039 0 diode
R46040 N46039 N46040 10
D46040 N46040 0 diode
R46041 N46040 N46041 10
D46041 N46041 0 diode
R46042 N46041 N46042 10
D46042 N46042 0 diode
R46043 N46042 N46043 10
D46043 N46043 0 diode
R46044 N46043 N46044 10
D46044 N46044 0 diode
R46045 N46044 N46045 10
D46045 N46045 0 diode
R46046 N46045 N46046 10
D46046 N46046 0 diode
R46047 N46046 N46047 10
D46047 N46047 0 diode
R46048 N46047 N46048 10
D46048 N46048 0 diode
R46049 N46048 N46049 10
D46049 N46049 0 diode
R46050 N46049 N46050 10
D46050 N46050 0 diode
R46051 N46050 N46051 10
D46051 N46051 0 diode
R46052 N46051 N46052 10
D46052 N46052 0 diode
R46053 N46052 N46053 10
D46053 N46053 0 diode
R46054 N46053 N46054 10
D46054 N46054 0 diode
R46055 N46054 N46055 10
D46055 N46055 0 diode
R46056 N46055 N46056 10
D46056 N46056 0 diode
R46057 N46056 N46057 10
D46057 N46057 0 diode
R46058 N46057 N46058 10
D46058 N46058 0 diode
R46059 N46058 N46059 10
D46059 N46059 0 diode
R46060 N46059 N46060 10
D46060 N46060 0 diode
R46061 N46060 N46061 10
D46061 N46061 0 diode
R46062 N46061 N46062 10
D46062 N46062 0 diode
R46063 N46062 N46063 10
D46063 N46063 0 diode
R46064 N46063 N46064 10
D46064 N46064 0 diode
R46065 N46064 N46065 10
D46065 N46065 0 diode
R46066 N46065 N46066 10
D46066 N46066 0 diode
R46067 N46066 N46067 10
D46067 N46067 0 diode
R46068 N46067 N46068 10
D46068 N46068 0 diode
R46069 N46068 N46069 10
D46069 N46069 0 diode
R46070 N46069 N46070 10
D46070 N46070 0 diode
R46071 N46070 N46071 10
D46071 N46071 0 diode
R46072 N46071 N46072 10
D46072 N46072 0 diode
R46073 N46072 N46073 10
D46073 N46073 0 diode
R46074 N46073 N46074 10
D46074 N46074 0 diode
R46075 N46074 N46075 10
D46075 N46075 0 diode
R46076 N46075 N46076 10
D46076 N46076 0 diode
R46077 N46076 N46077 10
D46077 N46077 0 diode
R46078 N46077 N46078 10
D46078 N46078 0 diode
R46079 N46078 N46079 10
D46079 N46079 0 diode
R46080 N46079 N46080 10
D46080 N46080 0 diode
R46081 N46080 N46081 10
D46081 N46081 0 diode
R46082 N46081 N46082 10
D46082 N46082 0 diode
R46083 N46082 N46083 10
D46083 N46083 0 diode
R46084 N46083 N46084 10
D46084 N46084 0 diode
R46085 N46084 N46085 10
D46085 N46085 0 diode
R46086 N46085 N46086 10
D46086 N46086 0 diode
R46087 N46086 N46087 10
D46087 N46087 0 diode
R46088 N46087 N46088 10
D46088 N46088 0 diode
R46089 N46088 N46089 10
D46089 N46089 0 diode
R46090 N46089 N46090 10
D46090 N46090 0 diode
R46091 N46090 N46091 10
D46091 N46091 0 diode
R46092 N46091 N46092 10
D46092 N46092 0 diode
R46093 N46092 N46093 10
D46093 N46093 0 diode
R46094 N46093 N46094 10
D46094 N46094 0 diode
R46095 N46094 N46095 10
D46095 N46095 0 diode
R46096 N46095 N46096 10
D46096 N46096 0 diode
R46097 N46096 N46097 10
D46097 N46097 0 diode
R46098 N46097 N46098 10
D46098 N46098 0 diode
R46099 N46098 N46099 10
D46099 N46099 0 diode
R46100 N46099 N46100 10
D46100 N46100 0 diode
R46101 N46100 N46101 10
D46101 N46101 0 diode
R46102 N46101 N46102 10
D46102 N46102 0 diode
R46103 N46102 N46103 10
D46103 N46103 0 diode
R46104 N46103 N46104 10
D46104 N46104 0 diode
R46105 N46104 N46105 10
D46105 N46105 0 diode
R46106 N46105 N46106 10
D46106 N46106 0 diode
R46107 N46106 N46107 10
D46107 N46107 0 diode
R46108 N46107 N46108 10
D46108 N46108 0 diode
R46109 N46108 N46109 10
D46109 N46109 0 diode
R46110 N46109 N46110 10
D46110 N46110 0 diode
R46111 N46110 N46111 10
D46111 N46111 0 diode
R46112 N46111 N46112 10
D46112 N46112 0 diode
R46113 N46112 N46113 10
D46113 N46113 0 diode
R46114 N46113 N46114 10
D46114 N46114 0 diode
R46115 N46114 N46115 10
D46115 N46115 0 diode
R46116 N46115 N46116 10
D46116 N46116 0 diode
R46117 N46116 N46117 10
D46117 N46117 0 diode
R46118 N46117 N46118 10
D46118 N46118 0 diode
R46119 N46118 N46119 10
D46119 N46119 0 diode
R46120 N46119 N46120 10
D46120 N46120 0 diode
R46121 N46120 N46121 10
D46121 N46121 0 diode
R46122 N46121 N46122 10
D46122 N46122 0 diode
R46123 N46122 N46123 10
D46123 N46123 0 diode
R46124 N46123 N46124 10
D46124 N46124 0 diode
R46125 N46124 N46125 10
D46125 N46125 0 diode
R46126 N46125 N46126 10
D46126 N46126 0 diode
R46127 N46126 N46127 10
D46127 N46127 0 diode
R46128 N46127 N46128 10
D46128 N46128 0 diode
R46129 N46128 N46129 10
D46129 N46129 0 diode
R46130 N46129 N46130 10
D46130 N46130 0 diode
R46131 N46130 N46131 10
D46131 N46131 0 diode
R46132 N46131 N46132 10
D46132 N46132 0 diode
R46133 N46132 N46133 10
D46133 N46133 0 diode
R46134 N46133 N46134 10
D46134 N46134 0 diode
R46135 N46134 N46135 10
D46135 N46135 0 diode
R46136 N46135 N46136 10
D46136 N46136 0 diode
R46137 N46136 N46137 10
D46137 N46137 0 diode
R46138 N46137 N46138 10
D46138 N46138 0 diode
R46139 N46138 N46139 10
D46139 N46139 0 diode
R46140 N46139 N46140 10
D46140 N46140 0 diode
R46141 N46140 N46141 10
D46141 N46141 0 diode
R46142 N46141 N46142 10
D46142 N46142 0 diode
R46143 N46142 N46143 10
D46143 N46143 0 diode
R46144 N46143 N46144 10
D46144 N46144 0 diode
R46145 N46144 N46145 10
D46145 N46145 0 diode
R46146 N46145 N46146 10
D46146 N46146 0 diode
R46147 N46146 N46147 10
D46147 N46147 0 diode
R46148 N46147 N46148 10
D46148 N46148 0 diode
R46149 N46148 N46149 10
D46149 N46149 0 diode
R46150 N46149 N46150 10
D46150 N46150 0 diode
R46151 N46150 N46151 10
D46151 N46151 0 diode
R46152 N46151 N46152 10
D46152 N46152 0 diode
R46153 N46152 N46153 10
D46153 N46153 0 diode
R46154 N46153 N46154 10
D46154 N46154 0 diode
R46155 N46154 N46155 10
D46155 N46155 0 diode
R46156 N46155 N46156 10
D46156 N46156 0 diode
R46157 N46156 N46157 10
D46157 N46157 0 diode
R46158 N46157 N46158 10
D46158 N46158 0 diode
R46159 N46158 N46159 10
D46159 N46159 0 diode
R46160 N46159 N46160 10
D46160 N46160 0 diode
R46161 N46160 N46161 10
D46161 N46161 0 diode
R46162 N46161 N46162 10
D46162 N46162 0 diode
R46163 N46162 N46163 10
D46163 N46163 0 diode
R46164 N46163 N46164 10
D46164 N46164 0 diode
R46165 N46164 N46165 10
D46165 N46165 0 diode
R46166 N46165 N46166 10
D46166 N46166 0 diode
R46167 N46166 N46167 10
D46167 N46167 0 diode
R46168 N46167 N46168 10
D46168 N46168 0 diode
R46169 N46168 N46169 10
D46169 N46169 0 diode
R46170 N46169 N46170 10
D46170 N46170 0 diode
R46171 N46170 N46171 10
D46171 N46171 0 diode
R46172 N46171 N46172 10
D46172 N46172 0 diode
R46173 N46172 N46173 10
D46173 N46173 0 diode
R46174 N46173 N46174 10
D46174 N46174 0 diode
R46175 N46174 N46175 10
D46175 N46175 0 diode
R46176 N46175 N46176 10
D46176 N46176 0 diode
R46177 N46176 N46177 10
D46177 N46177 0 diode
R46178 N46177 N46178 10
D46178 N46178 0 diode
R46179 N46178 N46179 10
D46179 N46179 0 diode
R46180 N46179 N46180 10
D46180 N46180 0 diode
R46181 N46180 N46181 10
D46181 N46181 0 diode
R46182 N46181 N46182 10
D46182 N46182 0 diode
R46183 N46182 N46183 10
D46183 N46183 0 diode
R46184 N46183 N46184 10
D46184 N46184 0 diode
R46185 N46184 N46185 10
D46185 N46185 0 diode
R46186 N46185 N46186 10
D46186 N46186 0 diode
R46187 N46186 N46187 10
D46187 N46187 0 diode
R46188 N46187 N46188 10
D46188 N46188 0 diode
R46189 N46188 N46189 10
D46189 N46189 0 diode
R46190 N46189 N46190 10
D46190 N46190 0 diode
R46191 N46190 N46191 10
D46191 N46191 0 diode
R46192 N46191 N46192 10
D46192 N46192 0 diode
R46193 N46192 N46193 10
D46193 N46193 0 diode
R46194 N46193 N46194 10
D46194 N46194 0 diode
R46195 N46194 N46195 10
D46195 N46195 0 diode
R46196 N46195 N46196 10
D46196 N46196 0 diode
R46197 N46196 N46197 10
D46197 N46197 0 diode
R46198 N46197 N46198 10
D46198 N46198 0 diode
R46199 N46198 N46199 10
D46199 N46199 0 diode
R46200 N46199 N46200 10
D46200 N46200 0 diode
R46201 N46200 N46201 10
D46201 N46201 0 diode
R46202 N46201 N46202 10
D46202 N46202 0 diode
R46203 N46202 N46203 10
D46203 N46203 0 diode
R46204 N46203 N46204 10
D46204 N46204 0 diode
R46205 N46204 N46205 10
D46205 N46205 0 diode
R46206 N46205 N46206 10
D46206 N46206 0 diode
R46207 N46206 N46207 10
D46207 N46207 0 diode
R46208 N46207 N46208 10
D46208 N46208 0 diode
R46209 N46208 N46209 10
D46209 N46209 0 diode
R46210 N46209 N46210 10
D46210 N46210 0 diode
R46211 N46210 N46211 10
D46211 N46211 0 diode
R46212 N46211 N46212 10
D46212 N46212 0 diode
R46213 N46212 N46213 10
D46213 N46213 0 diode
R46214 N46213 N46214 10
D46214 N46214 0 diode
R46215 N46214 N46215 10
D46215 N46215 0 diode
R46216 N46215 N46216 10
D46216 N46216 0 diode
R46217 N46216 N46217 10
D46217 N46217 0 diode
R46218 N46217 N46218 10
D46218 N46218 0 diode
R46219 N46218 N46219 10
D46219 N46219 0 diode
R46220 N46219 N46220 10
D46220 N46220 0 diode
R46221 N46220 N46221 10
D46221 N46221 0 diode
R46222 N46221 N46222 10
D46222 N46222 0 diode
R46223 N46222 N46223 10
D46223 N46223 0 diode
R46224 N46223 N46224 10
D46224 N46224 0 diode
R46225 N46224 N46225 10
D46225 N46225 0 diode
R46226 N46225 N46226 10
D46226 N46226 0 diode
R46227 N46226 N46227 10
D46227 N46227 0 diode
R46228 N46227 N46228 10
D46228 N46228 0 diode
R46229 N46228 N46229 10
D46229 N46229 0 diode
R46230 N46229 N46230 10
D46230 N46230 0 diode
R46231 N46230 N46231 10
D46231 N46231 0 diode
R46232 N46231 N46232 10
D46232 N46232 0 diode
R46233 N46232 N46233 10
D46233 N46233 0 diode
R46234 N46233 N46234 10
D46234 N46234 0 diode
R46235 N46234 N46235 10
D46235 N46235 0 diode
R46236 N46235 N46236 10
D46236 N46236 0 diode
R46237 N46236 N46237 10
D46237 N46237 0 diode
R46238 N46237 N46238 10
D46238 N46238 0 diode
R46239 N46238 N46239 10
D46239 N46239 0 diode
R46240 N46239 N46240 10
D46240 N46240 0 diode
R46241 N46240 N46241 10
D46241 N46241 0 diode
R46242 N46241 N46242 10
D46242 N46242 0 diode
R46243 N46242 N46243 10
D46243 N46243 0 diode
R46244 N46243 N46244 10
D46244 N46244 0 diode
R46245 N46244 N46245 10
D46245 N46245 0 diode
R46246 N46245 N46246 10
D46246 N46246 0 diode
R46247 N46246 N46247 10
D46247 N46247 0 diode
R46248 N46247 N46248 10
D46248 N46248 0 diode
R46249 N46248 N46249 10
D46249 N46249 0 diode
R46250 N46249 N46250 10
D46250 N46250 0 diode
R46251 N46250 N46251 10
D46251 N46251 0 diode
R46252 N46251 N46252 10
D46252 N46252 0 diode
R46253 N46252 N46253 10
D46253 N46253 0 diode
R46254 N46253 N46254 10
D46254 N46254 0 diode
R46255 N46254 N46255 10
D46255 N46255 0 diode
R46256 N46255 N46256 10
D46256 N46256 0 diode
R46257 N46256 N46257 10
D46257 N46257 0 diode
R46258 N46257 N46258 10
D46258 N46258 0 diode
R46259 N46258 N46259 10
D46259 N46259 0 diode
R46260 N46259 N46260 10
D46260 N46260 0 diode
R46261 N46260 N46261 10
D46261 N46261 0 diode
R46262 N46261 N46262 10
D46262 N46262 0 diode
R46263 N46262 N46263 10
D46263 N46263 0 diode
R46264 N46263 N46264 10
D46264 N46264 0 diode
R46265 N46264 N46265 10
D46265 N46265 0 diode
R46266 N46265 N46266 10
D46266 N46266 0 diode
R46267 N46266 N46267 10
D46267 N46267 0 diode
R46268 N46267 N46268 10
D46268 N46268 0 diode
R46269 N46268 N46269 10
D46269 N46269 0 diode
R46270 N46269 N46270 10
D46270 N46270 0 diode
R46271 N46270 N46271 10
D46271 N46271 0 diode
R46272 N46271 N46272 10
D46272 N46272 0 diode
R46273 N46272 N46273 10
D46273 N46273 0 diode
R46274 N46273 N46274 10
D46274 N46274 0 diode
R46275 N46274 N46275 10
D46275 N46275 0 diode
R46276 N46275 N46276 10
D46276 N46276 0 diode
R46277 N46276 N46277 10
D46277 N46277 0 diode
R46278 N46277 N46278 10
D46278 N46278 0 diode
R46279 N46278 N46279 10
D46279 N46279 0 diode
R46280 N46279 N46280 10
D46280 N46280 0 diode
R46281 N46280 N46281 10
D46281 N46281 0 diode
R46282 N46281 N46282 10
D46282 N46282 0 diode
R46283 N46282 N46283 10
D46283 N46283 0 diode
R46284 N46283 N46284 10
D46284 N46284 0 diode
R46285 N46284 N46285 10
D46285 N46285 0 diode
R46286 N46285 N46286 10
D46286 N46286 0 diode
R46287 N46286 N46287 10
D46287 N46287 0 diode
R46288 N46287 N46288 10
D46288 N46288 0 diode
R46289 N46288 N46289 10
D46289 N46289 0 diode
R46290 N46289 N46290 10
D46290 N46290 0 diode
R46291 N46290 N46291 10
D46291 N46291 0 diode
R46292 N46291 N46292 10
D46292 N46292 0 diode
R46293 N46292 N46293 10
D46293 N46293 0 diode
R46294 N46293 N46294 10
D46294 N46294 0 diode
R46295 N46294 N46295 10
D46295 N46295 0 diode
R46296 N46295 N46296 10
D46296 N46296 0 diode
R46297 N46296 N46297 10
D46297 N46297 0 diode
R46298 N46297 N46298 10
D46298 N46298 0 diode
R46299 N46298 N46299 10
D46299 N46299 0 diode
R46300 N46299 N46300 10
D46300 N46300 0 diode
R46301 N46300 N46301 10
D46301 N46301 0 diode
R46302 N46301 N46302 10
D46302 N46302 0 diode
R46303 N46302 N46303 10
D46303 N46303 0 diode
R46304 N46303 N46304 10
D46304 N46304 0 diode
R46305 N46304 N46305 10
D46305 N46305 0 diode
R46306 N46305 N46306 10
D46306 N46306 0 diode
R46307 N46306 N46307 10
D46307 N46307 0 diode
R46308 N46307 N46308 10
D46308 N46308 0 diode
R46309 N46308 N46309 10
D46309 N46309 0 diode
R46310 N46309 N46310 10
D46310 N46310 0 diode
R46311 N46310 N46311 10
D46311 N46311 0 diode
R46312 N46311 N46312 10
D46312 N46312 0 diode
R46313 N46312 N46313 10
D46313 N46313 0 diode
R46314 N46313 N46314 10
D46314 N46314 0 diode
R46315 N46314 N46315 10
D46315 N46315 0 diode
R46316 N46315 N46316 10
D46316 N46316 0 diode
R46317 N46316 N46317 10
D46317 N46317 0 diode
R46318 N46317 N46318 10
D46318 N46318 0 diode
R46319 N46318 N46319 10
D46319 N46319 0 diode
R46320 N46319 N46320 10
D46320 N46320 0 diode
R46321 N46320 N46321 10
D46321 N46321 0 diode
R46322 N46321 N46322 10
D46322 N46322 0 diode
R46323 N46322 N46323 10
D46323 N46323 0 diode
R46324 N46323 N46324 10
D46324 N46324 0 diode
R46325 N46324 N46325 10
D46325 N46325 0 diode
R46326 N46325 N46326 10
D46326 N46326 0 diode
R46327 N46326 N46327 10
D46327 N46327 0 diode
R46328 N46327 N46328 10
D46328 N46328 0 diode
R46329 N46328 N46329 10
D46329 N46329 0 diode
R46330 N46329 N46330 10
D46330 N46330 0 diode
R46331 N46330 N46331 10
D46331 N46331 0 diode
R46332 N46331 N46332 10
D46332 N46332 0 diode
R46333 N46332 N46333 10
D46333 N46333 0 diode
R46334 N46333 N46334 10
D46334 N46334 0 diode
R46335 N46334 N46335 10
D46335 N46335 0 diode
R46336 N46335 N46336 10
D46336 N46336 0 diode
R46337 N46336 N46337 10
D46337 N46337 0 diode
R46338 N46337 N46338 10
D46338 N46338 0 diode
R46339 N46338 N46339 10
D46339 N46339 0 diode
R46340 N46339 N46340 10
D46340 N46340 0 diode
R46341 N46340 N46341 10
D46341 N46341 0 diode
R46342 N46341 N46342 10
D46342 N46342 0 diode
R46343 N46342 N46343 10
D46343 N46343 0 diode
R46344 N46343 N46344 10
D46344 N46344 0 diode
R46345 N46344 N46345 10
D46345 N46345 0 diode
R46346 N46345 N46346 10
D46346 N46346 0 diode
R46347 N46346 N46347 10
D46347 N46347 0 diode
R46348 N46347 N46348 10
D46348 N46348 0 diode
R46349 N46348 N46349 10
D46349 N46349 0 diode
R46350 N46349 N46350 10
D46350 N46350 0 diode
R46351 N46350 N46351 10
D46351 N46351 0 diode
R46352 N46351 N46352 10
D46352 N46352 0 diode
R46353 N46352 N46353 10
D46353 N46353 0 diode
R46354 N46353 N46354 10
D46354 N46354 0 diode
R46355 N46354 N46355 10
D46355 N46355 0 diode
R46356 N46355 N46356 10
D46356 N46356 0 diode
R46357 N46356 N46357 10
D46357 N46357 0 diode
R46358 N46357 N46358 10
D46358 N46358 0 diode
R46359 N46358 N46359 10
D46359 N46359 0 diode
R46360 N46359 N46360 10
D46360 N46360 0 diode
R46361 N46360 N46361 10
D46361 N46361 0 diode
R46362 N46361 N46362 10
D46362 N46362 0 diode
R46363 N46362 N46363 10
D46363 N46363 0 diode
R46364 N46363 N46364 10
D46364 N46364 0 diode
R46365 N46364 N46365 10
D46365 N46365 0 diode
R46366 N46365 N46366 10
D46366 N46366 0 diode
R46367 N46366 N46367 10
D46367 N46367 0 diode
R46368 N46367 N46368 10
D46368 N46368 0 diode
R46369 N46368 N46369 10
D46369 N46369 0 diode
R46370 N46369 N46370 10
D46370 N46370 0 diode
R46371 N46370 N46371 10
D46371 N46371 0 diode
R46372 N46371 N46372 10
D46372 N46372 0 diode
R46373 N46372 N46373 10
D46373 N46373 0 diode
R46374 N46373 N46374 10
D46374 N46374 0 diode
R46375 N46374 N46375 10
D46375 N46375 0 diode
R46376 N46375 N46376 10
D46376 N46376 0 diode
R46377 N46376 N46377 10
D46377 N46377 0 diode
R46378 N46377 N46378 10
D46378 N46378 0 diode
R46379 N46378 N46379 10
D46379 N46379 0 diode
R46380 N46379 N46380 10
D46380 N46380 0 diode
R46381 N46380 N46381 10
D46381 N46381 0 diode
R46382 N46381 N46382 10
D46382 N46382 0 diode
R46383 N46382 N46383 10
D46383 N46383 0 diode
R46384 N46383 N46384 10
D46384 N46384 0 diode
R46385 N46384 N46385 10
D46385 N46385 0 diode
R46386 N46385 N46386 10
D46386 N46386 0 diode
R46387 N46386 N46387 10
D46387 N46387 0 diode
R46388 N46387 N46388 10
D46388 N46388 0 diode
R46389 N46388 N46389 10
D46389 N46389 0 diode
R46390 N46389 N46390 10
D46390 N46390 0 diode
R46391 N46390 N46391 10
D46391 N46391 0 diode
R46392 N46391 N46392 10
D46392 N46392 0 diode
R46393 N46392 N46393 10
D46393 N46393 0 diode
R46394 N46393 N46394 10
D46394 N46394 0 diode
R46395 N46394 N46395 10
D46395 N46395 0 diode
R46396 N46395 N46396 10
D46396 N46396 0 diode
R46397 N46396 N46397 10
D46397 N46397 0 diode
R46398 N46397 N46398 10
D46398 N46398 0 diode
R46399 N46398 N46399 10
D46399 N46399 0 diode
R46400 N46399 N46400 10
D46400 N46400 0 diode
R46401 N46400 N46401 10
D46401 N46401 0 diode
R46402 N46401 N46402 10
D46402 N46402 0 diode
R46403 N46402 N46403 10
D46403 N46403 0 diode
R46404 N46403 N46404 10
D46404 N46404 0 diode
R46405 N46404 N46405 10
D46405 N46405 0 diode
R46406 N46405 N46406 10
D46406 N46406 0 diode
R46407 N46406 N46407 10
D46407 N46407 0 diode
R46408 N46407 N46408 10
D46408 N46408 0 diode
R46409 N46408 N46409 10
D46409 N46409 0 diode
R46410 N46409 N46410 10
D46410 N46410 0 diode
R46411 N46410 N46411 10
D46411 N46411 0 diode
R46412 N46411 N46412 10
D46412 N46412 0 diode
R46413 N46412 N46413 10
D46413 N46413 0 diode
R46414 N46413 N46414 10
D46414 N46414 0 diode
R46415 N46414 N46415 10
D46415 N46415 0 diode
R46416 N46415 N46416 10
D46416 N46416 0 diode
R46417 N46416 N46417 10
D46417 N46417 0 diode
R46418 N46417 N46418 10
D46418 N46418 0 diode
R46419 N46418 N46419 10
D46419 N46419 0 diode
R46420 N46419 N46420 10
D46420 N46420 0 diode
R46421 N46420 N46421 10
D46421 N46421 0 diode
R46422 N46421 N46422 10
D46422 N46422 0 diode
R46423 N46422 N46423 10
D46423 N46423 0 diode
R46424 N46423 N46424 10
D46424 N46424 0 diode
R46425 N46424 N46425 10
D46425 N46425 0 diode
R46426 N46425 N46426 10
D46426 N46426 0 diode
R46427 N46426 N46427 10
D46427 N46427 0 diode
R46428 N46427 N46428 10
D46428 N46428 0 diode
R46429 N46428 N46429 10
D46429 N46429 0 diode
R46430 N46429 N46430 10
D46430 N46430 0 diode
R46431 N46430 N46431 10
D46431 N46431 0 diode
R46432 N46431 N46432 10
D46432 N46432 0 diode
R46433 N46432 N46433 10
D46433 N46433 0 diode
R46434 N46433 N46434 10
D46434 N46434 0 diode
R46435 N46434 N46435 10
D46435 N46435 0 diode
R46436 N46435 N46436 10
D46436 N46436 0 diode
R46437 N46436 N46437 10
D46437 N46437 0 diode
R46438 N46437 N46438 10
D46438 N46438 0 diode
R46439 N46438 N46439 10
D46439 N46439 0 diode
R46440 N46439 N46440 10
D46440 N46440 0 diode
R46441 N46440 N46441 10
D46441 N46441 0 diode
R46442 N46441 N46442 10
D46442 N46442 0 diode
R46443 N46442 N46443 10
D46443 N46443 0 diode
R46444 N46443 N46444 10
D46444 N46444 0 diode
R46445 N46444 N46445 10
D46445 N46445 0 diode
R46446 N46445 N46446 10
D46446 N46446 0 diode
R46447 N46446 N46447 10
D46447 N46447 0 diode
R46448 N46447 N46448 10
D46448 N46448 0 diode
R46449 N46448 N46449 10
D46449 N46449 0 diode
R46450 N46449 N46450 10
D46450 N46450 0 diode
R46451 N46450 N46451 10
D46451 N46451 0 diode
R46452 N46451 N46452 10
D46452 N46452 0 diode
R46453 N46452 N46453 10
D46453 N46453 0 diode
R46454 N46453 N46454 10
D46454 N46454 0 diode
R46455 N46454 N46455 10
D46455 N46455 0 diode
R46456 N46455 N46456 10
D46456 N46456 0 diode
R46457 N46456 N46457 10
D46457 N46457 0 diode
R46458 N46457 N46458 10
D46458 N46458 0 diode
R46459 N46458 N46459 10
D46459 N46459 0 diode
R46460 N46459 N46460 10
D46460 N46460 0 diode
R46461 N46460 N46461 10
D46461 N46461 0 diode
R46462 N46461 N46462 10
D46462 N46462 0 diode
R46463 N46462 N46463 10
D46463 N46463 0 diode
R46464 N46463 N46464 10
D46464 N46464 0 diode
R46465 N46464 N46465 10
D46465 N46465 0 diode
R46466 N46465 N46466 10
D46466 N46466 0 diode
R46467 N46466 N46467 10
D46467 N46467 0 diode
R46468 N46467 N46468 10
D46468 N46468 0 diode
R46469 N46468 N46469 10
D46469 N46469 0 diode
R46470 N46469 N46470 10
D46470 N46470 0 diode
R46471 N46470 N46471 10
D46471 N46471 0 diode
R46472 N46471 N46472 10
D46472 N46472 0 diode
R46473 N46472 N46473 10
D46473 N46473 0 diode
R46474 N46473 N46474 10
D46474 N46474 0 diode
R46475 N46474 N46475 10
D46475 N46475 0 diode
R46476 N46475 N46476 10
D46476 N46476 0 diode
R46477 N46476 N46477 10
D46477 N46477 0 diode
R46478 N46477 N46478 10
D46478 N46478 0 diode
R46479 N46478 N46479 10
D46479 N46479 0 diode
R46480 N46479 N46480 10
D46480 N46480 0 diode
R46481 N46480 N46481 10
D46481 N46481 0 diode
R46482 N46481 N46482 10
D46482 N46482 0 diode
R46483 N46482 N46483 10
D46483 N46483 0 diode
R46484 N46483 N46484 10
D46484 N46484 0 diode
R46485 N46484 N46485 10
D46485 N46485 0 diode
R46486 N46485 N46486 10
D46486 N46486 0 diode
R46487 N46486 N46487 10
D46487 N46487 0 diode
R46488 N46487 N46488 10
D46488 N46488 0 diode
R46489 N46488 N46489 10
D46489 N46489 0 diode
R46490 N46489 N46490 10
D46490 N46490 0 diode
R46491 N46490 N46491 10
D46491 N46491 0 diode
R46492 N46491 N46492 10
D46492 N46492 0 diode
R46493 N46492 N46493 10
D46493 N46493 0 diode
R46494 N46493 N46494 10
D46494 N46494 0 diode
R46495 N46494 N46495 10
D46495 N46495 0 diode
R46496 N46495 N46496 10
D46496 N46496 0 diode
R46497 N46496 N46497 10
D46497 N46497 0 diode
R46498 N46497 N46498 10
D46498 N46498 0 diode
R46499 N46498 N46499 10
D46499 N46499 0 diode
R46500 N46499 N46500 10
D46500 N46500 0 diode
R46501 N46500 N46501 10
D46501 N46501 0 diode
R46502 N46501 N46502 10
D46502 N46502 0 diode
R46503 N46502 N46503 10
D46503 N46503 0 diode
R46504 N46503 N46504 10
D46504 N46504 0 diode
R46505 N46504 N46505 10
D46505 N46505 0 diode
R46506 N46505 N46506 10
D46506 N46506 0 diode
R46507 N46506 N46507 10
D46507 N46507 0 diode
R46508 N46507 N46508 10
D46508 N46508 0 diode
R46509 N46508 N46509 10
D46509 N46509 0 diode
R46510 N46509 N46510 10
D46510 N46510 0 diode
R46511 N46510 N46511 10
D46511 N46511 0 diode
R46512 N46511 N46512 10
D46512 N46512 0 diode
R46513 N46512 N46513 10
D46513 N46513 0 diode
R46514 N46513 N46514 10
D46514 N46514 0 diode
R46515 N46514 N46515 10
D46515 N46515 0 diode
R46516 N46515 N46516 10
D46516 N46516 0 diode
R46517 N46516 N46517 10
D46517 N46517 0 diode
R46518 N46517 N46518 10
D46518 N46518 0 diode
R46519 N46518 N46519 10
D46519 N46519 0 diode
R46520 N46519 N46520 10
D46520 N46520 0 diode
R46521 N46520 N46521 10
D46521 N46521 0 diode
R46522 N46521 N46522 10
D46522 N46522 0 diode
R46523 N46522 N46523 10
D46523 N46523 0 diode
R46524 N46523 N46524 10
D46524 N46524 0 diode
R46525 N46524 N46525 10
D46525 N46525 0 diode
R46526 N46525 N46526 10
D46526 N46526 0 diode
R46527 N46526 N46527 10
D46527 N46527 0 diode
R46528 N46527 N46528 10
D46528 N46528 0 diode
R46529 N46528 N46529 10
D46529 N46529 0 diode
R46530 N46529 N46530 10
D46530 N46530 0 diode
R46531 N46530 N46531 10
D46531 N46531 0 diode
R46532 N46531 N46532 10
D46532 N46532 0 diode
R46533 N46532 N46533 10
D46533 N46533 0 diode
R46534 N46533 N46534 10
D46534 N46534 0 diode
R46535 N46534 N46535 10
D46535 N46535 0 diode
R46536 N46535 N46536 10
D46536 N46536 0 diode
R46537 N46536 N46537 10
D46537 N46537 0 diode
R46538 N46537 N46538 10
D46538 N46538 0 diode
R46539 N46538 N46539 10
D46539 N46539 0 diode
R46540 N46539 N46540 10
D46540 N46540 0 diode
R46541 N46540 N46541 10
D46541 N46541 0 diode
R46542 N46541 N46542 10
D46542 N46542 0 diode
R46543 N46542 N46543 10
D46543 N46543 0 diode
R46544 N46543 N46544 10
D46544 N46544 0 diode
R46545 N46544 N46545 10
D46545 N46545 0 diode
R46546 N46545 N46546 10
D46546 N46546 0 diode
R46547 N46546 N46547 10
D46547 N46547 0 diode
R46548 N46547 N46548 10
D46548 N46548 0 diode
R46549 N46548 N46549 10
D46549 N46549 0 diode
R46550 N46549 N46550 10
D46550 N46550 0 diode
R46551 N46550 N46551 10
D46551 N46551 0 diode
R46552 N46551 N46552 10
D46552 N46552 0 diode
R46553 N46552 N46553 10
D46553 N46553 0 diode
R46554 N46553 N46554 10
D46554 N46554 0 diode
R46555 N46554 N46555 10
D46555 N46555 0 diode
R46556 N46555 N46556 10
D46556 N46556 0 diode
R46557 N46556 N46557 10
D46557 N46557 0 diode
R46558 N46557 N46558 10
D46558 N46558 0 diode
R46559 N46558 N46559 10
D46559 N46559 0 diode
R46560 N46559 N46560 10
D46560 N46560 0 diode
R46561 N46560 N46561 10
D46561 N46561 0 diode
R46562 N46561 N46562 10
D46562 N46562 0 diode
R46563 N46562 N46563 10
D46563 N46563 0 diode
R46564 N46563 N46564 10
D46564 N46564 0 diode
R46565 N46564 N46565 10
D46565 N46565 0 diode
R46566 N46565 N46566 10
D46566 N46566 0 diode
R46567 N46566 N46567 10
D46567 N46567 0 diode
R46568 N46567 N46568 10
D46568 N46568 0 diode
R46569 N46568 N46569 10
D46569 N46569 0 diode
R46570 N46569 N46570 10
D46570 N46570 0 diode
R46571 N46570 N46571 10
D46571 N46571 0 diode
R46572 N46571 N46572 10
D46572 N46572 0 diode
R46573 N46572 N46573 10
D46573 N46573 0 diode
R46574 N46573 N46574 10
D46574 N46574 0 diode
R46575 N46574 N46575 10
D46575 N46575 0 diode
R46576 N46575 N46576 10
D46576 N46576 0 diode
R46577 N46576 N46577 10
D46577 N46577 0 diode
R46578 N46577 N46578 10
D46578 N46578 0 diode
R46579 N46578 N46579 10
D46579 N46579 0 diode
R46580 N46579 N46580 10
D46580 N46580 0 diode
R46581 N46580 N46581 10
D46581 N46581 0 diode
R46582 N46581 N46582 10
D46582 N46582 0 diode
R46583 N46582 N46583 10
D46583 N46583 0 diode
R46584 N46583 N46584 10
D46584 N46584 0 diode
R46585 N46584 N46585 10
D46585 N46585 0 diode
R46586 N46585 N46586 10
D46586 N46586 0 diode
R46587 N46586 N46587 10
D46587 N46587 0 diode
R46588 N46587 N46588 10
D46588 N46588 0 diode
R46589 N46588 N46589 10
D46589 N46589 0 diode
R46590 N46589 N46590 10
D46590 N46590 0 diode
R46591 N46590 N46591 10
D46591 N46591 0 diode
R46592 N46591 N46592 10
D46592 N46592 0 diode
R46593 N46592 N46593 10
D46593 N46593 0 diode
R46594 N46593 N46594 10
D46594 N46594 0 diode
R46595 N46594 N46595 10
D46595 N46595 0 diode
R46596 N46595 N46596 10
D46596 N46596 0 diode
R46597 N46596 N46597 10
D46597 N46597 0 diode
R46598 N46597 N46598 10
D46598 N46598 0 diode
R46599 N46598 N46599 10
D46599 N46599 0 diode
R46600 N46599 N46600 10
D46600 N46600 0 diode
R46601 N46600 N46601 10
D46601 N46601 0 diode
R46602 N46601 N46602 10
D46602 N46602 0 diode
R46603 N46602 N46603 10
D46603 N46603 0 diode
R46604 N46603 N46604 10
D46604 N46604 0 diode
R46605 N46604 N46605 10
D46605 N46605 0 diode
R46606 N46605 N46606 10
D46606 N46606 0 diode
R46607 N46606 N46607 10
D46607 N46607 0 diode
R46608 N46607 N46608 10
D46608 N46608 0 diode
R46609 N46608 N46609 10
D46609 N46609 0 diode
R46610 N46609 N46610 10
D46610 N46610 0 diode
R46611 N46610 N46611 10
D46611 N46611 0 diode
R46612 N46611 N46612 10
D46612 N46612 0 diode
R46613 N46612 N46613 10
D46613 N46613 0 diode
R46614 N46613 N46614 10
D46614 N46614 0 diode
R46615 N46614 N46615 10
D46615 N46615 0 diode
R46616 N46615 N46616 10
D46616 N46616 0 diode
R46617 N46616 N46617 10
D46617 N46617 0 diode
R46618 N46617 N46618 10
D46618 N46618 0 diode
R46619 N46618 N46619 10
D46619 N46619 0 diode
R46620 N46619 N46620 10
D46620 N46620 0 diode
R46621 N46620 N46621 10
D46621 N46621 0 diode
R46622 N46621 N46622 10
D46622 N46622 0 diode
R46623 N46622 N46623 10
D46623 N46623 0 diode
R46624 N46623 N46624 10
D46624 N46624 0 diode
R46625 N46624 N46625 10
D46625 N46625 0 diode
R46626 N46625 N46626 10
D46626 N46626 0 diode
R46627 N46626 N46627 10
D46627 N46627 0 diode
R46628 N46627 N46628 10
D46628 N46628 0 diode
R46629 N46628 N46629 10
D46629 N46629 0 diode
R46630 N46629 N46630 10
D46630 N46630 0 diode
R46631 N46630 N46631 10
D46631 N46631 0 diode
R46632 N46631 N46632 10
D46632 N46632 0 diode
R46633 N46632 N46633 10
D46633 N46633 0 diode
R46634 N46633 N46634 10
D46634 N46634 0 diode
R46635 N46634 N46635 10
D46635 N46635 0 diode
R46636 N46635 N46636 10
D46636 N46636 0 diode
R46637 N46636 N46637 10
D46637 N46637 0 diode
R46638 N46637 N46638 10
D46638 N46638 0 diode
R46639 N46638 N46639 10
D46639 N46639 0 diode
R46640 N46639 N46640 10
D46640 N46640 0 diode
R46641 N46640 N46641 10
D46641 N46641 0 diode
R46642 N46641 N46642 10
D46642 N46642 0 diode
R46643 N46642 N46643 10
D46643 N46643 0 diode
R46644 N46643 N46644 10
D46644 N46644 0 diode
R46645 N46644 N46645 10
D46645 N46645 0 diode
R46646 N46645 N46646 10
D46646 N46646 0 diode
R46647 N46646 N46647 10
D46647 N46647 0 diode
R46648 N46647 N46648 10
D46648 N46648 0 diode
R46649 N46648 N46649 10
D46649 N46649 0 diode
R46650 N46649 N46650 10
D46650 N46650 0 diode
R46651 N46650 N46651 10
D46651 N46651 0 diode
R46652 N46651 N46652 10
D46652 N46652 0 diode
R46653 N46652 N46653 10
D46653 N46653 0 diode
R46654 N46653 N46654 10
D46654 N46654 0 diode
R46655 N46654 N46655 10
D46655 N46655 0 diode
R46656 N46655 N46656 10
D46656 N46656 0 diode
R46657 N46656 N46657 10
D46657 N46657 0 diode
R46658 N46657 N46658 10
D46658 N46658 0 diode
R46659 N46658 N46659 10
D46659 N46659 0 diode
R46660 N46659 N46660 10
D46660 N46660 0 diode
R46661 N46660 N46661 10
D46661 N46661 0 diode
R46662 N46661 N46662 10
D46662 N46662 0 diode
R46663 N46662 N46663 10
D46663 N46663 0 diode
R46664 N46663 N46664 10
D46664 N46664 0 diode
R46665 N46664 N46665 10
D46665 N46665 0 diode
R46666 N46665 N46666 10
D46666 N46666 0 diode
R46667 N46666 N46667 10
D46667 N46667 0 diode
R46668 N46667 N46668 10
D46668 N46668 0 diode
R46669 N46668 N46669 10
D46669 N46669 0 diode
R46670 N46669 N46670 10
D46670 N46670 0 diode
R46671 N46670 N46671 10
D46671 N46671 0 diode
R46672 N46671 N46672 10
D46672 N46672 0 diode
R46673 N46672 N46673 10
D46673 N46673 0 diode
R46674 N46673 N46674 10
D46674 N46674 0 diode
R46675 N46674 N46675 10
D46675 N46675 0 diode
R46676 N46675 N46676 10
D46676 N46676 0 diode
R46677 N46676 N46677 10
D46677 N46677 0 diode
R46678 N46677 N46678 10
D46678 N46678 0 diode
R46679 N46678 N46679 10
D46679 N46679 0 diode
R46680 N46679 N46680 10
D46680 N46680 0 diode
R46681 N46680 N46681 10
D46681 N46681 0 diode
R46682 N46681 N46682 10
D46682 N46682 0 diode
R46683 N46682 N46683 10
D46683 N46683 0 diode
R46684 N46683 N46684 10
D46684 N46684 0 diode
R46685 N46684 N46685 10
D46685 N46685 0 diode
R46686 N46685 N46686 10
D46686 N46686 0 diode
R46687 N46686 N46687 10
D46687 N46687 0 diode
R46688 N46687 N46688 10
D46688 N46688 0 diode
R46689 N46688 N46689 10
D46689 N46689 0 diode
R46690 N46689 N46690 10
D46690 N46690 0 diode
R46691 N46690 N46691 10
D46691 N46691 0 diode
R46692 N46691 N46692 10
D46692 N46692 0 diode
R46693 N46692 N46693 10
D46693 N46693 0 diode
R46694 N46693 N46694 10
D46694 N46694 0 diode
R46695 N46694 N46695 10
D46695 N46695 0 diode
R46696 N46695 N46696 10
D46696 N46696 0 diode
R46697 N46696 N46697 10
D46697 N46697 0 diode
R46698 N46697 N46698 10
D46698 N46698 0 diode
R46699 N46698 N46699 10
D46699 N46699 0 diode
R46700 N46699 N46700 10
D46700 N46700 0 diode
R46701 N46700 N46701 10
D46701 N46701 0 diode
R46702 N46701 N46702 10
D46702 N46702 0 diode
R46703 N46702 N46703 10
D46703 N46703 0 diode
R46704 N46703 N46704 10
D46704 N46704 0 diode
R46705 N46704 N46705 10
D46705 N46705 0 diode
R46706 N46705 N46706 10
D46706 N46706 0 diode
R46707 N46706 N46707 10
D46707 N46707 0 diode
R46708 N46707 N46708 10
D46708 N46708 0 diode
R46709 N46708 N46709 10
D46709 N46709 0 diode
R46710 N46709 N46710 10
D46710 N46710 0 diode
R46711 N46710 N46711 10
D46711 N46711 0 diode
R46712 N46711 N46712 10
D46712 N46712 0 diode
R46713 N46712 N46713 10
D46713 N46713 0 diode
R46714 N46713 N46714 10
D46714 N46714 0 diode
R46715 N46714 N46715 10
D46715 N46715 0 diode
R46716 N46715 N46716 10
D46716 N46716 0 diode
R46717 N46716 N46717 10
D46717 N46717 0 diode
R46718 N46717 N46718 10
D46718 N46718 0 diode
R46719 N46718 N46719 10
D46719 N46719 0 diode
R46720 N46719 N46720 10
D46720 N46720 0 diode
R46721 N46720 N46721 10
D46721 N46721 0 diode
R46722 N46721 N46722 10
D46722 N46722 0 diode
R46723 N46722 N46723 10
D46723 N46723 0 diode
R46724 N46723 N46724 10
D46724 N46724 0 diode
R46725 N46724 N46725 10
D46725 N46725 0 diode
R46726 N46725 N46726 10
D46726 N46726 0 diode
R46727 N46726 N46727 10
D46727 N46727 0 diode
R46728 N46727 N46728 10
D46728 N46728 0 diode
R46729 N46728 N46729 10
D46729 N46729 0 diode
R46730 N46729 N46730 10
D46730 N46730 0 diode
R46731 N46730 N46731 10
D46731 N46731 0 diode
R46732 N46731 N46732 10
D46732 N46732 0 diode
R46733 N46732 N46733 10
D46733 N46733 0 diode
R46734 N46733 N46734 10
D46734 N46734 0 diode
R46735 N46734 N46735 10
D46735 N46735 0 diode
R46736 N46735 N46736 10
D46736 N46736 0 diode
R46737 N46736 N46737 10
D46737 N46737 0 diode
R46738 N46737 N46738 10
D46738 N46738 0 diode
R46739 N46738 N46739 10
D46739 N46739 0 diode
R46740 N46739 N46740 10
D46740 N46740 0 diode
R46741 N46740 N46741 10
D46741 N46741 0 diode
R46742 N46741 N46742 10
D46742 N46742 0 diode
R46743 N46742 N46743 10
D46743 N46743 0 diode
R46744 N46743 N46744 10
D46744 N46744 0 diode
R46745 N46744 N46745 10
D46745 N46745 0 diode
R46746 N46745 N46746 10
D46746 N46746 0 diode
R46747 N46746 N46747 10
D46747 N46747 0 diode
R46748 N46747 N46748 10
D46748 N46748 0 diode
R46749 N46748 N46749 10
D46749 N46749 0 diode
R46750 N46749 N46750 10
D46750 N46750 0 diode
R46751 N46750 N46751 10
D46751 N46751 0 diode
R46752 N46751 N46752 10
D46752 N46752 0 diode
R46753 N46752 N46753 10
D46753 N46753 0 diode
R46754 N46753 N46754 10
D46754 N46754 0 diode
R46755 N46754 N46755 10
D46755 N46755 0 diode
R46756 N46755 N46756 10
D46756 N46756 0 diode
R46757 N46756 N46757 10
D46757 N46757 0 diode
R46758 N46757 N46758 10
D46758 N46758 0 diode
R46759 N46758 N46759 10
D46759 N46759 0 diode
R46760 N46759 N46760 10
D46760 N46760 0 diode
R46761 N46760 N46761 10
D46761 N46761 0 diode
R46762 N46761 N46762 10
D46762 N46762 0 diode
R46763 N46762 N46763 10
D46763 N46763 0 diode
R46764 N46763 N46764 10
D46764 N46764 0 diode
R46765 N46764 N46765 10
D46765 N46765 0 diode
R46766 N46765 N46766 10
D46766 N46766 0 diode
R46767 N46766 N46767 10
D46767 N46767 0 diode
R46768 N46767 N46768 10
D46768 N46768 0 diode
R46769 N46768 N46769 10
D46769 N46769 0 diode
R46770 N46769 N46770 10
D46770 N46770 0 diode
R46771 N46770 N46771 10
D46771 N46771 0 diode
R46772 N46771 N46772 10
D46772 N46772 0 diode
R46773 N46772 N46773 10
D46773 N46773 0 diode
R46774 N46773 N46774 10
D46774 N46774 0 diode
R46775 N46774 N46775 10
D46775 N46775 0 diode
R46776 N46775 N46776 10
D46776 N46776 0 diode
R46777 N46776 N46777 10
D46777 N46777 0 diode
R46778 N46777 N46778 10
D46778 N46778 0 diode
R46779 N46778 N46779 10
D46779 N46779 0 diode
R46780 N46779 N46780 10
D46780 N46780 0 diode
R46781 N46780 N46781 10
D46781 N46781 0 diode
R46782 N46781 N46782 10
D46782 N46782 0 diode
R46783 N46782 N46783 10
D46783 N46783 0 diode
R46784 N46783 N46784 10
D46784 N46784 0 diode
R46785 N46784 N46785 10
D46785 N46785 0 diode
R46786 N46785 N46786 10
D46786 N46786 0 diode
R46787 N46786 N46787 10
D46787 N46787 0 diode
R46788 N46787 N46788 10
D46788 N46788 0 diode
R46789 N46788 N46789 10
D46789 N46789 0 diode
R46790 N46789 N46790 10
D46790 N46790 0 diode
R46791 N46790 N46791 10
D46791 N46791 0 diode
R46792 N46791 N46792 10
D46792 N46792 0 diode
R46793 N46792 N46793 10
D46793 N46793 0 diode
R46794 N46793 N46794 10
D46794 N46794 0 diode
R46795 N46794 N46795 10
D46795 N46795 0 diode
R46796 N46795 N46796 10
D46796 N46796 0 diode
R46797 N46796 N46797 10
D46797 N46797 0 diode
R46798 N46797 N46798 10
D46798 N46798 0 diode
R46799 N46798 N46799 10
D46799 N46799 0 diode
R46800 N46799 N46800 10
D46800 N46800 0 diode
R46801 N46800 N46801 10
D46801 N46801 0 diode
R46802 N46801 N46802 10
D46802 N46802 0 diode
R46803 N46802 N46803 10
D46803 N46803 0 diode
R46804 N46803 N46804 10
D46804 N46804 0 diode
R46805 N46804 N46805 10
D46805 N46805 0 diode
R46806 N46805 N46806 10
D46806 N46806 0 diode
R46807 N46806 N46807 10
D46807 N46807 0 diode
R46808 N46807 N46808 10
D46808 N46808 0 diode
R46809 N46808 N46809 10
D46809 N46809 0 diode
R46810 N46809 N46810 10
D46810 N46810 0 diode
R46811 N46810 N46811 10
D46811 N46811 0 diode
R46812 N46811 N46812 10
D46812 N46812 0 diode
R46813 N46812 N46813 10
D46813 N46813 0 diode
R46814 N46813 N46814 10
D46814 N46814 0 diode
R46815 N46814 N46815 10
D46815 N46815 0 diode
R46816 N46815 N46816 10
D46816 N46816 0 diode
R46817 N46816 N46817 10
D46817 N46817 0 diode
R46818 N46817 N46818 10
D46818 N46818 0 diode
R46819 N46818 N46819 10
D46819 N46819 0 diode
R46820 N46819 N46820 10
D46820 N46820 0 diode
R46821 N46820 N46821 10
D46821 N46821 0 diode
R46822 N46821 N46822 10
D46822 N46822 0 diode
R46823 N46822 N46823 10
D46823 N46823 0 diode
R46824 N46823 N46824 10
D46824 N46824 0 diode
R46825 N46824 N46825 10
D46825 N46825 0 diode
R46826 N46825 N46826 10
D46826 N46826 0 diode
R46827 N46826 N46827 10
D46827 N46827 0 diode
R46828 N46827 N46828 10
D46828 N46828 0 diode
R46829 N46828 N46829 10
D46829 N46829 0 diode
R46830 N46829 N46830 10
D46830 N46830 0 diode
R46831 N46830 N46831 10
D46831 N46831 0 diode
R46832 N46831 N46832 10
D46832 N46832 0 diode
R46833 N46832 N46833 10
D46833 N46833 0 diode
R46834 N46833 N46834 10
D46834 N46834 0 diode
R46835 N46834 N46835 10
D46835 N46835 0 diode
R46836 N46835 N46836 10
D46836 N46836 0 diode
R46837 N46836 N46837 10
D46837 N46837 0 diode
R46838 N46837 N46838 10
D46838 N46838 0 diode
R46839 N46838 N46839 10
D46839 N46839 0 diode
R46840 N46839 N46840 10
D46840 N46840 0 diode
R46841 N46840 N46841 10
D46841 N46841 0 diode
R46842 N46841 N46842 10
D46842 N46842 0 diode
R46843 N46842 N46843 10
D46843 N46843 0 diode
R46844 N46843 N46844 10
D46844 N46844 0 diode
R46845 N46844 N46845 10
D46845 N46845 0 diode
R46846 N46845 N46846 10
D46846 N46846 0 diode
R46847 N46846 N46847 10
D46847 N46847 0 diode
R46848 N46847 N46848 10
D46848 N46848 0 diode
R46849 N46848 N46849 10
D46849 N46849 0 diode
R46850 N46849 N46850 10
D46850 N46850 0 diode
R46851 N46850 N46851 10
D46851 N46851 0 diode
R46852 N46851 N46852 10
D46852 N46852 0 diode
R46853 N46852 N46853 10
D46853 N46853 0 diode
R46854 N46853 N46854 10
D46854 N46854 0 diode
R46855 N46854 N46855 10
D46855 N46855 0 diode
R46856 N46855 N46856 10
D46856 N46856 0 diode
R46857 N46856 N46857 10
D46857 N46857 0 diode
R46858 N46857 N46858 10
D46858 N46858 0 diode
R46859 N46858 N46859 10
D46859 N46859 0 diode
R46860 N46859 N46860 10
D46860 N46860 0 diode
R46861 N46860 N46861 10
D46861 N46861 0 diode
R46862 N46861 N46862 10
D46862 N46862 0 diode
R46863 N46862 N46863 10
D46863 N46863 0 diode
R46864 N46863 N46864 10
D46864 N46864 0 diode
R46865 N46864 N46865 10
D46865 N46865 0 diode
R46866 N46865 N46866 10
D46866 N46866 0 diode
R46867 N46866 N46867 10
D46867 N46867 0 diode
R46868 N46867 N46868 10
D46868 N46868 0 diode
R46869 N46868 N46869 10
D46869 N46869 0 diode
R46870 N46869 N46870 10
D46870 N46870 0 diode
R46871 N46870 N46871 10
D46871 N46871 0 diode
R46872 N46871 N46872 10
D46872 N46872 0 diode
R46873 N46872 N46873 10
D46873 N46873 0 diode
R46874 N46873 N46874 10
D46874 N46874 0 diode
R46875 N46874 N46875 10
D46875 N46875 0 diode
R46876 N46875 N46876 10
D46876 N46876 0 diode
R46877 N46876 N46877 10
D46877 N46877 0 diode
R46878 N46877 N46878 10
D46878 N46878 0 diode
R46879 N46878 N46879 10
D46879 N46879 0 diode
R46880 N46879 N46880 10
D46880 N46880 0 diode
R46881 N46880 N46881 10
D46881 N46881 0 diode
R46882 N46881 N46882 10
D46882 N46882 0 diode
R46883 N46882 N46883 10
D46883 N46883 0 diode
R46884 N46883 N46884 10
D46884 N46884 0 diode
R46885 N46884 N46885 10
D46885 N46885 0 diode
R46886 N46885 N46886 10
D46886 N46886 0 diode
R46887 N46886 N46887 10
D46887 N46887 0 diode
R46888 N46887 N46888 10
D46888 N46888 0 diode
R46889 N46888 N46889 10
D46889 N46889 0 diode
R46890 N46889 N46890 10
D46890 N46890 0 diode
R46891 N46890 N46891 10
D46891 N46891 0 diode
R46892 N46891 N46892 10
D46892 N46892 0 diode
R46893 N46892 N46893 10
D46893 N46893 0 diode
R46894 N46893 N46894 10
D46894 N46894 0 diode
R46895 N46894 N46895 10
D46895 N46895 0 diode
R46896 N46895 N46896 10
D46896 N46896 0 diode
R46897 N46896 N46897 10
D46897 N46897 0 diode
R46898 N46897 N46898 10
D46898 N46898 0 diode
R46899 N46898 N46899 10
D46899 N46899 0 diode
R46900 N46899 N46900 10
D46900 N46900 0 diode
R46901 N46900 N46901 10
D46901 N46901 0 diode
R46902 N46901 N46902 10
D46902 N46902 0 diode
R46903 N46902 N46903 10
D46903 N46903 0 diode
R46904 N46903 N46904 10
D46904 N46904 0 diode
R46905 N46904 N46905 10
D46905 N46905 0 diode
R46906 N46905 N46906 10
D46906 N46906 0 diode
R46907 N46906 N46907 10
D46907 N46907 0 diode
R46908 N46907 N46908 10
D46908 N46908 0 diode
R46909 N46908 N46909 10
D46909 N46909 0 diode
R46910 N46909 N46910 10
D46910 N46910 0 diode
R46911 N46910 N46911 10
D46911 N46911 0 diode
R46912 N46911 N46912 10
D46912 N46912 0 diode
R46913 N46912 N46913 10
D46913 N46913 0 diode
R46914 N46913 N46914 10
D46914 N46914 0 diode
R46915 N46914 N46915 10
D46915 N46915 0 diode
R46916 N46915 N46916 10
D46916 N46916 0 diode
R46917 N46916 N46917 10
D46917 N46917 0 diode
R46918 N46917 N46918 10
D46918 N46918 0 diode
R46919 N46918 N46919 10
D46919 N46919 0 diode
R46920 N46919 N46920 10
D46920 N46920 0 diode
R46921 N46920 N46921 10
D46921 N46921 0 diode
R46922 N46921 N46922 10
D46922 N46922 0 diode
R46923 N46922 N46923 10
D46923 N46923 0 diode
R46924 N46923 N46924 10
D46924 N46924 0 diode
R46925 N46924 N46925 10
D46925 N46925 0 diode
R46926 N46925 N46926 10
D46926 N46926 0 diode
R46927 N46926 N46927 10
D46927 N46927 0 diode
R46928 N46927 N46928 10
D46928 N46928 0 diode
R46929 N46928 N46929 10
D46929 N46929 0 diode
R46930 N46929 N46930 10
D46930 N46930 0 diode
R46931 N46930 N46931 10
D46931 N46931 0 diode
R46932 N46931 N46932 10
D46932 N46932 0 diode
R46933 N46932 N46933 10
D46933 N46933 0 diode
R46934 N46933 N46934 10
D46934 N46934 0 diode
R46935 N46934 N46935 10
D46935 N46935 0 diode
R46936 N46935 N46936 10
D46936 N46936 0 diode
R46937 N46936 N46937 10
D46937 N46937 0 diode
R46938 N46937 N46938 10
D46938 N46938 0 diode
R46939 N46938 N46939 10
D46939 N46939 0 diode
R46940 N46939 N46940 10
D46940 N46940 0 diode
R46941 N46940 N46941 10
D46941 N46941 0 diode
R46942 N46941 N46942 10
D46942 N46942 0 diode
R46943 N46942 N46943 10
D46943 N46943 0 diode
R46944 N46943 N46944 10
D46944 N46944 0 diode
R46945 N46944 N46945 10
D46945 N46945 0 diode
R46946 N46945 N46946 10
D46946 N46946 0 diode
R46947 N46946 N46947 10
D46947 N46947 0 diode
R46948 N46947 N46948 10
D46948 N46948 0 diode
R46949 N46948 N46949 10
D46949 N46949 0 diode
R46950 N46949 N46950 10
D46950 N46950 0 diode
R46951 N46950 N46951 10
D46951 N46951 0 diode
R46952 N46951 N46952 10
D46952 N46952 0 diode
R46953 N46952 N46953 10
D46953 N46953 0 diode
R46954 N46953 N46954 10
D46954 N46954 0 diode
R46955 N46954 N46955 10
D46955 N46955 0 diode
R46956 N46955 N46956 10
D46956 N46956 0 diode
R46957 N46956 N46957 10
D46957 N46957 0 diode
R46958 N46957 N46958 10
D46958 N46958 0 diode
R46959 N46958 N46959 10
D46959 N46959 0 diode
R46960 N46959 N46960 10
D46960 N46960 0 diode
R46961 N46960 N46961 10
D46961 N46961 0 diode
R46962 N46961 N46962 10
D46962 N46962 0 diode
R46963 N46962 N46963 10
D46963 N46963 0 diode
R46964 N46963 N46964 10
D46964 N46964 0 diode
R46965 N46964 N46965 10
D46965 N46965 0 diode
R46966 N46965 N46966 10
D46966 N46966 0 diode
R46967 N46966 N46967 10
D46967 N46967 0 diode
R46968 N46967 N46968 10
D46968 N46968 0 diode
R46969 N46968 N46969 10
D46969 N46969 0 diode
R46970 N46969 N46970 10
D46970 N46970 0 diode
R46971 N46970 N46971 10
D46971 N46971 0 diode
R46972 N46971 N46972 10
D46972 N46972 0 diode
R46973 N46972 N46973 10
D46973 N46973 0 diode
R46974 N46973 N46974 10
D46974 N46974 0 diode
R46975 N46974 N46975 10
D46975 N46975 0 diode
R46976 N46975 N46976 10
D46976 N46976 0 diode
R46977 N46976 N46977 10
D46977 N46977 0 diode
R46978 N46977 N46978 10
D46978 N46978 0 diode
R46979 N46978 N46979 10
D46979 N46979 0 diode
R46980 N46979 N46980 10
D46980 N46980 0 diode
R46981 N46980 N46981 10
D46981 N46981 0 diode
R46982 N46981 N46982 10
D46982 N46982 0 diode
R46983 N46982 N46983 10
D46983 N46983 0 diode
R46984 N46983 N46984 10
D46984 N46984 0 diode
R46985 N46984 N46985 10
D46985 N46985 0 diode
R46986 N46985 N46986 10
D46986 N46986 0 diode
R46987 N46986 N46987 10
D46987 N46987 0 diode
R46988 N46987 N46988 10
D46988 N46988 0 diode
R46989 N46988 N46989 10
D46989 N46989 0 diode
R46990 N46989 N46990 10
D46990 N46990 0 diode
R46991 N46990 N46991 10
D46991 N46991 0 diode
R46992 N46991 N46992 10
D46992 N46992 0 diode
R46993 N46992 N46993 10
D46993 N46993 0 diode
R46994 N46993 N46994 10
D46994 N46994 0 diode
R46995 N46994 N46995 10
D46995 N46995 0 diode
R46996 N46995 N46996 10
D46996 N46996 0 diode
R46997 N46996 N46997 10
D46997 N46997 0 diode
R46998 N46997 N46998 10
D46998 N46998 0 diode
R46999 N46998 N46999 10
D46999 N46999 0 diode
R47000 N46999 N47000 10
D47000 N47000 0 diode
R47001 N47000 N47001 10
D47001 N47001 0 diode
R47002 N47001 N47002 10
D47002 N47002 0 diode
R47003 N47002 N47003 10
D47003 N47003 0 diode
R47004 N47003 N47004 10
D47004 N47004 0 diode
R47005 N47004 N47005 10
D47005 N47005 0 diode
R47006 N47005 N47006 10
D47006 N47006 0 diode
R47007 N47006 N47007 10
D47007 N47007 0 diode
R47008 N47007 N47008 10
D47008 N47008 0 diode
R47009 N47008 N47009 10
D47009 N47009 0 diode
R47010 N47009 N47010 10
D47010 N47010 0 diode
R47011 N47010 N47011 10
D47011 N47011 0 diode
R47012 N47011 N47012 10
D47012 N47012 0 diode
R47013 N47012 N47013 10
D47013 N47013 0 diode
R47014 N47013 N47014 10
D47014 N47014 0 diode
R47015 N47014 N47015 10
D47015 N47015 0 diode
R47016 N47015 N47016 10
D47016 N47016 0 diode
R47017 N47016 N47017 10
D47017 N47017 0 diode
R47018 N47017 N47018 10
D47018 N47018 0 diode
R47019 N47018 N47019 10
D47019 N47019 0 diode
R47020 N47019 N47020 10
D47020 N47020 0 diode
R47021 N47020 N47021 10
D47021 N47021 0 diode
R47022 N47021 N47022 10
D47022 N47022 0 diode
R47023 N47022 N47023 10
D47023 N47023 0 diode
R47024 N47023 N47024 10
D47024 N47024 0 diode
R47025 N47024 N47025 10
D47025 N47025 0 diode
R47026 N47025 N47026 10
D47026 N47026 0 diode
R47027 N47026 N47027 10
D47027 N47027 0 diode
R47028 N47027 N47028 10
D47028 N47028 0 diode
R47029 N47028 N47029 10
D47029 N47029 0 diode
R47030 N47029 N47030 10
D47030 N47030 0 diode
R47031 N47030 N47031 10
D47031 N47031 0 diode
R47032 N47031 N47032 10
D47032 N47032 0 diode
R47033 N47032 N47033 10
D47033 N47033 0 diode
R47034 N47033 N47034 10
D47034 N47034 0 diode
R47035 N47034 N47035 10
D47035 N47035 0 diode
R47036 N47035 N47036 10
D47036 N47036 0 diode
R47037 N47036 N47037 10
D47037 N47037 0 diode
R47038 N47037 N47038 10
D47038 N47038 0 diode
R47039 N47038 N47039 10
D47039 N47039 0 diode
R47040 N47039 N47040 10
D47040 N47040 0 diode
R47041 N47040 N47041 10
D47041 N47041 0 diode
R47042 N47041 N47042 10
D47042 N47042 0 diode
R47043 N47042 N47043 10
D47043 N47043 0 diode
R47044 N47043 N47044 10
D47044 N47044 0 diode
R47045 N47044 N47045 10
D47045 N47045 0 diode
R47046 N47045 N47046 10
D47046 N47046 0 diode
R47047 N47046 N47047 10
D47047 N47047 0 diode
R47048 N47047 N47048 10
D47048 N47048 0 diode
R47049 N47048 N47049 10
D47049 N47049 0 diode
R47050 N47049 N47050 10
D47050 N47050 0 diode
R47051 N47050 N47051 10
D47051 N47051 0 diode
R47052 N47051 N47052 10
D47052 N47052 0 diode
R47053 N47052 N47053 10
D47053 N47053 0 diode
R47054 N47053 N47054 10
D47054 N47054 0 diode
R47055 N47054 N47055 10
D47055 N47055 0 diode
R47056 N47055 N47056 10
D47056 N47056 0 diode
R47057 N47056 N47057 10
D47057 N47057 0 diode
R47058 N47057 N47058 10
D47058 N47058 0 diode
R47059 N47058 N47059 10
D47059 N47059 0 diode
R47060 N47059 N47060 10
D47060 N47060 0 diode
R47061 N47060 N47061 10
D47061 N47061 0 diode
R47062 N47061 N47062 10
D47062 N47062 0 diode
R47063 N47062 N47063 10
D47063 N47063 0 diode
R47064 N47063 N47064 10
D47064 N47064 0 diode
R47065 N47064 N47065 10
D47065 N47065 0 diode
R47066 N47065 N47066 10
D47066 N47066 0 diode
R47067 N47066 N47067 10
D47067 N47067 0 diode
R47068 N47067 N47068 10
D47068 N47068 0 diode
R47069 N47068 N47069 10
D47069 N47069 0 diode
R47070 N47069 N47070 10
D47070 N47070 0 diode
R47071 N47070 N47071 10
D47071 N47071 0 diode
R47072 N47071 N47072 10
D47072 N47072 0 diode
R47073 N47072 N47073 10
D47073 N47073 0 diode
R47074 N47073 N47074 10
D47074 N47074 0 diode
R47075 N47074 N47075 10
D47075 N47075 0 diode
R47076 N47075 N47076 10
D47076 N47076 0 diode
R47077 N47076 N47077 10
D47077 N47077 0 diode
R47078 N47077 N47078 10
D47078 N47078 0 diode
R47079 N47078 N47079 10
D47079 N47079 0 diode
R47080 N47079 N47080 10
D47080 N47080 0 diode
R47081 N47080 N47081 10
D47081 N47081 0 diode
R47082 N47081 N47082 10
D47082 N47082 0 diode
R47083 N47082 N47083 10
D47083 N47083 0 diode
R47084 N47083 N47084 10
D47084 N47084 0 diode
R47085 N47084 N47085 10
D47085 N47085 0 diode
R47086 N47085 N47086 10
D47086 N47086 0 diode
R47087 N47086 N47087 10
D47087 N47087 0 diode
R47088 N47087 N47088 10
D47088 N47088 0 diode
R47089 N47088 N47089 10
D47089 N47089 0 diode
R47090 N47089 N47090 10
D47090 N47090 0 diode
R47091 N47090 N47091 10
D47091 N47091 0 diode
R47092 N47091 N47092 10
D47092 N47092 0 diode
R47093 N47092 N47093 10
D47093 N47093 0 diode
R47094 N47093 N47094 10
D47094 N47094 0 diode
R47095 N47094 N47095 10
D47095 N47095 0 diode
R47096 N47095 N47096 10
D47096 N47096 0 diode
R47097 N47096 N47097 10
D47097 N47097 0 diode
R47098 N47097 N47098 10
D47098 N47098 0 diode
R47099 N47098 N47099 10
D47099 N47099 0 diode
R47100 N47099 N47100 10
D47100 N47100 0 diode
R47101 N47100 N47101 10
D47101 N47101 0 diode
R47102 N47101 N47102 10
D47102 N47102 0 diode
R47103 N47102 N47103 10
D47103 N47103 0 diode
R47104 N47103 N47104 10
D47104 N47104 0 diode
R47105 N47104 N47105 10
D47105 N47105 0 diode
R47106 N47105 N47106 10
D47106 N47106 0 diode
R47107 N47106 N47107 10
D47107 N47107 0 diode
R47108 N47107 N47108 10
D47108 N47108 0 diode
R47109 N47108 N47109 10
D47109 N47109 0 diode
R47110 N47109 N47110 10
D47110 N47110 0 diode
R47111 N47110 N47111 10
D47111 N47111 0 diode
R47112 N47111 N47112 10
D47112 N47112 0 diode
R47113 N47112 N47113 10
D47113 N47113 0 diode
R47114 N47113 N47114 10
D47114 N47114 0 diode
R47115 N47114 N47115 10
D47115 N47115 0 diode
R47116 N47115 N47116 10
D47116 N47116 0 diode
R47117 N47116 N47117 10
D47117 N47117 0 diode
R47118 N47117 N47118 10
D47118 N47118 0 diode
R47119 N47118 N47119 10
D47119 N47119 0 diode
R47120 N47119 N47120 10
D47120 N47120 0 diode
R47121 N47120 N47121 10
D47121 N47121 0 diode
R47122 N47121 N47122 10
D47122 N47122 0 diode
R47123 N47122 N47123 10
D47123 N47123 0 diode
R47124 N47123 N47124 10
D47124 N47124 0 diode
R47125 N47124 N47125 10
D47125 N47125 0 diode
R47126 N47125 N47126 10
D47126 N47126 0 diode
R47127 N47126 N47127 10
D47127 N47127 0 diode
R47128 N47127 N47128 10
D47128 N47128 0 diode
R47129 N47128 N47129 10
D47129 N47129 0 diode
R47130 N47129 N47130 10
D47130 N47130 0 diode
R47131 N47130 N47131 10
D47131 N47131 0 diode
R47132 N47131 N47132 10
D47132 N47132 0 diode
R47133 N47132 N47133 10
D47133 N47133 0 diode
R47134 N47133 N47134 10
D47134 N47134 0 diode
R47135 N47134 N47135 10
D47135 N47135 0 diode
R47136 N47135 N47136 10
D47136 N47136 0 diode
R47137 N47136 N47137 10
D47137 N47137 0 diode
R47138 N47137 N47138 10
D47138 N47138 0 diode
R47139 N47138 N47139 10
D47139 N47139 0 diode
R47140 N47139 N47140 10
D47140 N47140 0 diode
R47141 N47140 N47141 10
D47141 N47141 0 diode
R47142 N47141 N47142 10
D47142 N47142 0 diode
R47143 N47142 N47143 10
D47143 N47143 0 diode
R47144 N47143 N47144 10
D47144 N47144 0 diode
R47145 N47144 N47145 10
D47145 N47145 0 diode
R47146 N47145 N47146 10
D47146 N47146 0 diode
R47147 N47146 N47147 10
D47147 N47147 0 diode
R47148 N47147 N47148 10
D47148 N47148 0 diode
R47149 N47148 N47149 10
D47149 N47149 0 diode
R47150 N47149 N47150 10
D47150 N47150 0 diode
R47151 N47150 N47151 10
D47151 N47151 0 diode
R47152 N47151 N47152 10
D47152 N47152 0 diode
R47153 N47152 N47153 10
D47153 N47153 0 diode
R47154 N47153 N47154 10
D47154 N47154 0 diode
R47155 N47154 N47155 10
D47155 N47155 0 diode
R47156 N47155 N47156 10
D47156 N47156 0 diode
R47157 N47156 N47157 10
D47157 N47157 0 diode
R47158 N47157 N47158 10
D47158 N47158 0 diode
R47159 N47158 N47159 10
D47159 N47159 0 diode
R47160 N47159 N47160 10
D47160 N47160 0 diode
R47161 N47160 N47161 10
D47161 N47161 0 diode
R47162 N47161 N47162 10
D47162 N47162 0 diode
R47163 N47162 N47163 10
D47163 N47163 0 diode
R47164 N47163 N47164 10
D47164 N47164 0 diode
R47165 N47164 N47165 10
D47165 N47165 0 diode
R47166 N47165 N47166 10
D47166 N47166 0 diode
R47167 N47166 N47167 10
D47167 N47167 0 diode
R47168 N47167 N47168 10
D47168 N47168 0 diode
R47169 N47168 N47169 10
D47169 N47169 0 diode
R47170 N47169 N47170 10
D47170 N47170 0 diode
R47171 N47170 N47171 10
D47171 N47171 0 diode
R47172 N47171 N47172 10
D47172 N47172 0 diode
R47173 N47172 N47173 10
D47173 N47173 0 diode
R47174 N47173 N47174 10
D47174 N47174 0 diode
R47175 N47174 N47175 10
D47175 N47175 0 diode
R47176 N47175 N47176 10
D47176 N47176 0 diode
R47177 N47176 N47177 10
D47177 N47177 0 diode
R47178 N47177 N47178 10
D47178 N47178 0 diode
R47179 N47178 N47179 10
D47179 N47179 0 diode
R47180 N47179 N47180 10
D47180 N47180 0 diode
R47181 N47180 N47181 10
D47181 N47181 0 diode
R47182 N47181 N47182 10
D47182 N47182 0 diode
R47183 N47182 N47183 10
D47183 N47183 0 diode
R47184 N47183 N47184 10
D47184 N47184 0 diode
R47185 N47184 N47185 10
D47185 N47185 0 diode
R47186 N47185 N47186 10
D47186 N47186 0 diode
R47187 N47186 N47187 10
D47187 N47187 0 diode
R47188 N47187 N47188 10
D47188 N47188 0 diode
R47189 N47188 N47189 10
D47189 N47189 0 diode
R47190 N47189 N47190 10
D47190 N47190 0 diode
R47191 N47190 N47191 10
D47191 N47191 0 diode
R47192 N47191 N47192 10
D47192 N47192 0 diode
R47193 N47192 N47193 10
D47193 N47193 0 diode
R47194 N47193 N47194 10
D47194 N47194 0 diode
R47195 N47194 N47195 10
D47195 N47195 0 diode
R47196 N47195 N47196 10
D47196 N47196 0 diode
R47197 N47196 N47197 10
D47197 N47197 0 diode
R47198 N47197 N47198 10
D47198 N47198 0 diode
R47199 N47198 N47199 10
D47199 N47199 0 diode
R47200 N47199 N47200 10
D47200 N47200 0 diode
R47201 N47200 N47201 10
D47201 N47201 0 diode
R47202 N47201 N47202 10
D47202 N47202 0 diode
R47203 N47202 N47203 10
D47203 N47203 0 diode
R47204 N47203 N47204 10
D47204 N47204 0 diode
R47205 N47204 N47205 10
D47205 N47205 0 diode
R47206 N47205 N47206 10
D47206 N47206 0 diode
R47207 N47206 N47207 10
D47207 N47207 0 diode
R47208 N47207 N47208 10
D47208 N47208 0 diode
R47209 N47208 N47209 10
D47209 N47209 0 diode
R47210 N47209 N47210 10
D47210 N47210 0 diode
R47211 N47210 N47211 10
D47211 N47211 0 diode
R47212 N47211 N47212 10
D47212 N47212 0 diode
R47213 N47212 N47213 10
D47213 N47213 0 diode
R47214 N47213 N47214 10
D47214 N47214 0 diode
R47215 N47214 N47215 10
D47215 N47215 0 diode
R47216 N47215 N47216 10
D47216 N47216 0 diode
R47217 N47216 N47217 10
D47217 N47217 0 diode
R47218 N47217 N47218 10
D47218 N47218 0 diode
R47219 N47218 N47219 10
D47219 N47219 0 diode
R47220 N47219 N47220 10
D47220 N47220 0 diode
R47221 N47220 N47221 10
D47221 N47221 0 diode
R47222 N47221 N47222 10
D47222 N47222 0 diode
R47223 N47222 N47223 10
D47223 N47223 0 diode
R47224 N47223 N47224 10
D47224 N47224 0 diode
R47225 N47224 N47225 10
D47225 N47225 0 diode
R47226 N47225 N47226 10
D47226 N47226 0 diode
R47227 N47226 N47227 10
D47227 N47227 0 diode
R47228 N47227 N47228 10
D47228 N47228 0 diode
R47229 N47228 N47229 10
D47229 N47229 0 diode
R47230 N47229 N47230 10
D47230 N47230 0 diode
R47231 N47230 N47231 10
D47231 N47231 0 diode
R47232 N47231 N47232 10
D47232 N47232 0 diode
R47233 N47232 N47233 10
D47233 N47233 0 diode
R47234 N47233 N47234 10
D47234 N47234 0 diode
R47235 N47234 N47235 10
D47235 N47235 0 diode
R47236 N47235 N47236 10
D47236 N47236 0 diode
R47237 N47236 N47237 10
D47237 N47237 0 diode
R47238 N47237 N47238 10
D47238 N47238 0 diode
R47239 N47238 N47239 10
D47239 N47239 0 diode
R47240 N47239 N47240 10
D47240 N47240 0 diode
R47241 N47240 N47241 10
D47241 N47241 0 diode
R47242 N47241 N47242 10
D47242 N47242 0 diode
R47243 N47242 N47243 10
D47243 N47243 0 diode
R47244 N47243 N47244 10
D47244 N47244 0 diode
R47245 N47244 N47245 10
D47245 N47245 0 diode
R47246 N47245 N47246 10
D47246 N47246 0 diode
R47247 N47246 N47247 10
D47247 N47247 0 diode
R47248 N47247 N47248 10
D47248 N47248 0 diode
R47249 N47248 N47249 10
D47249 N47249 0 diode
R47250 N47249 N47250 10
D47250 N47250 0 diode
R47251 N47250 N47251 10
D47251 N47251 0 diode
R47252 N47251 N47252 10
D47252 N47252 0 diode
R47253 N47252 N47253 10
D47253 N47253 0 diode
R47254 N47253 N47254 10
D47254 N47254 0 diode
R47255 N47254 N47255 10
D47255 N47255 0 diode
R47256 N47255 N47256 10
D47256 N47256 0 diode
R47257 N47256 N47257 10
D47257 N47257 0 diode
R47258 N47257 N47258 10
D47258 N47258 0 diode
R47259 N47258 N47259 10
D47259 N47259 0 diode
R47260 N47259 N47260 10
D47260 N47260 0 diode
R47261 N47260 N47261 10
D47261 N47261 0 diode
R47262 N47261 N47262 10
D47262 N47262 0 diode
R47263 N47262 N47263 10
D47263 N47263 0 diode
R47264 N47263 N47264 10
D47264 N47264 0 diode
R47265 N47264 N47265 10
D47265 N47265 0 diode
R47266 N47265 N47266 10
D47266 N47266 0 diode
R47267 N47266 N47267 10
D47267 N47267 0 diode
R47268 N47267 N47268 10
D47268 N47268 0 diode
R47269 N47268 N47269 10
D47269 N47269 0 diode
R47270 N47269 N47270 10
D47270 N47270 0 diode
R47271 N47270 N47271 10
D47271 N47271 0 diode
R47272 N47271 N47272 10
D47272 N47272 0 diode
R47273 N47272 N47273 10
D47273 N47273 0 diode
R47274 N47273 N47274 10
D47274 N47274 0 diode
R47275 N47274 N47275 10
D47275 N47275 0 diode
R47276 N47275 N47276 10
D47276 N47276 0 diode
R47277 N47276 N47277 10
D47277 N47277 0 diode
R47278 N47277 N47278 10
D47278 N47278 0 diode
R47279 N47278 N47279 10
D47279 N47279 0 diode
R47280 N47279 N47280 10
D47280 N47280 0 diode
R47281 N47280 N47281 10
D47281 N47281 0 diode
R47282 N47281 N47282 10
D47282 N47282 0 diode
R47283 N47282 N47283 10
D47283 N47283 0 diode
R47284 N47283 N47284 10
D47284 N47284 0 diode
R47285 N47284 N47285 10
D47285 N47285 0 diode
R47286 N47285 N47286 10
D47286 N47286 0 diode
R47287 N47286 N47287 10
D47287 N47287 0 diode
R47288 N47287 N47288 10
D47288 N47288 0 diode
R47289 N47288 N47289 10
D47289 N47289 0 diode
R47290 N47289 N47290 10
D47290 N47290 0 diode
R47291 N47290 N47291 10
D47291 N47291 0 diode
R47292 N47291 N47292 10
D47292 N47292 0 diode
R47293 N47292 N47293 10
D47293 N47293 0 diode
R47294 N47293 N47294 10
D47294 N47294 0 diode
R47295 N47294 N47295 10
D47295 N47295 0 diode
R47296 N47295 N47296 10
D47296 N47296 0 diode
R47297 N47296 N47297 10
D47297 N47297 0 diode
R47298 N47297 N47298 10
D47298 N47298 0 diode
R47299 N47298 N47299 10
D47299 N47299 0 diode
R47300 N47299 N47300 10
D47300 N47300 0 diode
R47301 N47300 N47301 10
D47301 N47301 0 diode
R47302 N47301 N47302 10
D47302 N47302 0 diode
R47303 N47302 N47303 10
D47303 N47303 0 diode
R47304 N47303 N47304 10
D47304 N47304 0 diode
R47305 N47304 N47305 10
D47305 N47305 0 diode
R47306 N47305 N47306 10
D47306 N47306 0 diode
R47307 N47306 N47307 10
D47307 N47307 0 diode
R47308 N47307 N47308 10
D47308 N47308 0 diode
R47309 N47308 N47309 10
D47309 N47309 0 diode
R47310 N47309 N47310 10
D47310 N47310 0 diode
R47311 N47310 N47311 10
D47311 N47311 0 diode
R47312 N47311 N47312 10
D47312 N47312 0 diode
R47313 N47312 N47313 10
D47313 N47313 0 diode
R47314 N47313 N47314 10
D47314 N47314 0 diode
R47315 N47314 N47315 10
D47315 N47315 0 diode
R47316 N47315 N47316 10
D47316 N47316 0 diode
R47317 N47316 N47317 10
D47317 N47317 0 diode
R47318 N47317 N47318 10
D47318 N47318 0 diode
R47319 N47318 N47319 10
D47319 N47319 0 diode
R47320 N47319 N47320 10
D47320 N47320 0 diode
R47321 N47320 N47321 10
D47321 N47321 0 diode
R47322 N47321 N47322 10
D47322 N47322 0 diode
R47323 N47322 N47323 10
D47323 N47323 0 diode
R47324 N47323 N47324 10
D47324 N47324 0 diode
R47325 N47324 N47325 10
D47325 N47325 0 diode
R47326 N47325 N47326 10
D47326 N47326 0 diode
R47327 N47326 N47327 10
D47327 N47327 0 diode
R47328 N47327 N47328 10
D47328 N47328 0 diode
R47329 N47328 N47329 10
D47329 N47329 0 diode
R47330 N47329 N47330 10
D47330 N47330 0 diode
R47331 N47330 N47331 10
D47331 N47331 0 diode
R47332 N47331 N47332 10
D47332 N47332 0 diode
R47333 N47332 N47333 10
D47333 N47333 0 diode
R47334 N47333 N47334 10
D47334 N47334 0 diode
R47335 N47334 N47335 10
D47335 N47335 0 diode
R47336 N47335 N47336 10
D47336 N47336 0 diode
R47337 N47336 N47337 10
D47337 N47337 0 diode
R47338 N47337 N47338 10
D47338 N47338 0 diode
R47339 N47338 N47339 10
D47339 N47339 0 diode
R47340 N47339 N47340 10
D47340 N47340 0 diode
R47341 N47340 N47341 10
D47341 N47341 0 diode
R47342 N47341 N47342 10
D47342 N47342 0 diode
R47343 N47342 N47343 10
D47343 N47343 0 diode
R47344 N47343 N47344 10
D47344 N47344 0 diode
R47345 N47344 N47345 10
D47345 N47345 0 diode
R47346 N47345 N47346 10
D47346 N47346 0 diode
R47347 N47346 N47347 10
D47347 N47347 0 diode
R47348 N47347 N47348 10
D47348 N47348 0 diode
R47349 N47348 N47349 10
D47349 N47349 0 diode
R47350 N47349 N47350 10
D47350 N47350 0 diode
R47351 N47350 N47351 10
D47351 N47351 0 diode
R47352 N47351 N47352 10
D47352 N47352 0 diode
R47353 N47352 N47353 10
D47353 N47353 0 diode
R47354 N47353 N47354 10
D47354 N47354 0 diode
R47355 N47354 N47355 10
D47355 N47355 0 diode
R47356 N47355 N47356 10
D47356 N47356 0 diode
R47357 N47356 N47357 10
D47357 N47357 0 diode
R47358 N47357 N47358 10
D47358 N47358 0 diode
R47359 N47358 N47359 10
D47359 N47359 0 diode
R47360 N47359 N47360 10
D47360 N47360 0 diode
R47361 N47360 N47361 10
D47361 N47361 0 diode
R47362 N47361 N47362 10
D47362 N47362 0 diode
R47363 N47362 N47363 10
D47363 N47363 0 diode
R47364 N47363 N47364 10
D47364 N47364 0 diode
R47365 N47364 N47365 10
D47365 N47365 0 diode
R47366 N47365 N47366 10
D47366 N47366 0 diode
R47367 N47366 N47367 10
D47367 N47367 0 diode
R47368 N47367 N47368 10
D47368 N47368 0 diode
R47369 N47368 N47369 10
D47369 N47369 0 diode
R47370 N47369 N47370 10
D47370 N47370 0 diode
R47371 N47370 N47371 10
D47371 N47371 0 diode
R47372 N47371 N47372 10
D47372 N47372 0 diode
R47373 N47372 N47373 10
D47373 N47373 0 diode
R47374 N47373 N47374 10
D47374 N47374 0 diode
R47375 N47374 N47375 10
D47375 N47375 0 diode
R47376 N47375 N47376 10
D47376 N47376 0 diode
R47377 N47376 N47377 10
D47377 N47377 0 diode
R47378 N47377 N47378 10
D47378 N47378 0 diode
R47379 N47378 N47379 10
D47379 N47379 0 diode
R47380 N47379 N47380 10
D47380 N47380 0 diode
R47381 N47380 N47381 10
D47381 N47381 0 diode
R47382 N47381 N47382 10
D47382 N47382 0 diode
R47383 N47382 N47383 10
D47383 N47383 0 diode
R47384 N47383 N47384 10
D47384 N47384 0 diode
R47385 N47384 N47385 10
D47385 N47385 0 diode
R47386 N47385 N47386 10
D47386 N47386 0 diode
R47387 N47386 N47387 10
D47387 N47387 0 diode
R47388 N47387 N47388 10
D47388 N47388 0 diode
R47389 N47388 N47389 10
D47389 N47389 0 diode
R47390 N47389 N47390 10
D47390 N47390 0 diode
R47391 N47390 N47391 10
D47391 N47391 0 diode
R47392 N47391 N47392 10
D47392 N47392 0 diode
R47393 N47392 N47393 10
D47393 N47393 0 diode
R47394 N47393 N47394 10
D47394 N47394 0 diode
R47395 N47394 N47395 10
D47395 N47395 0 diode
R47396 N47395 N47396 10
D47396 N47396 0 diode
R47397 N47396 N47397 10
D47397 N47397 0 diode
R47398 N47397 N47398 10
D47398 N47398 0 diode
R47399 N47398 N47399 10
D47399 N47399 0 diode
R47400 N47399 N47400 10
D47400 N47400 0 diode
R47401 N47400 N47401 10
D47401 N47401 0 diode
R47402 N47401 N47402 10
D47402 N47402 0 diode
R47403 N47402 N47403 10
D47403 N47403 0 diode
R47404 N47403 N47404 10
D47404 N47404 0 diode
R47405 N47404 N47405 10
D47405 N47405 0 diode
R47406 N47405 N47406 10
D47406 N47406 0 diode
R47407 N47406 N47407 10
D47407 N47407 0 diode
R47408 N47407 N47408 10
D47408 N47408 0 diode
R47409 N47408 N47409 10
D47409 N47409 0 diode
R47410 N47409 N47410 10
D47410 N47410 0 diode
R47411 N47410 N47411 10
D47411 N47411 0 diode
R47412 N47411 N47412 10
D47412 N47412 0 diode
R47413 N47412 N47413 10
D47413 N47413 0 diode
R47414 N47413 N47414 10
D47414 N47414 0 diode
R47415 N47414 N47415 10
D47415 N47415 0 diode
R47416 N47415 N47416 10
D47416 N47416 0 diode
R47417 N47416 N47417 10
D47417 N47417 0 diode
R47418 N47417 N47418 10
D47418 N47418 0 diode
R47419 N47418 N47419 10
D47419 N47419 0 diode
R47420 N47419 N47420 10
D47420 N47420 0 diode
R47421 N47420 N47421 10
D47421 N47421 0 diode
R47422 N47421 N47422 10
D47422 N47422 0 diode
R47423 N47422 N47423 10
D47423 N47423 0 diode
R47424 N47423 N47424 10
D47424 N47424 0 diode
R47425 N47424 N47425 10
D47425 N47425 0 diode
R47426 N47425 N47426 10
D47426 N47426 0 diode
R47427 N47426 N47427 10
D47427 N47427 0 diode
R47428 N47427 N47428 10
D47428 N47428 0 diode
R47429 N47428 N47429 10
D47429 N47429 0 diode
R47430 N47429 N47430 10
D47430 N47430 0 diode
R47431 N47430 N47431 10
D47431 N47431 0 diode
R47432 N47431 N47432 10
D47432 N47432 0 diode
R47433 N47432 N47433 10
D47433 N47433 0 diode
R47434 N47433 N47434 10
D47434 N47434 0 diode
R47435 N47434 N47435 10
D47435 N47435 0 diode
R47436 N47435 N47436 10
D47436 N47436 0 diode
R47437 N47436 N47437 10
D47437 N47437 0 diode
R47438 N47437 N47438 10
D47438 N47438 0 diode
R47439 N47438 N47439 10
D47439 N47439 0 diode
R47440 N47439 N47440 10
D47440 N47440 0 diode
R47441 N47440 N47441 10
D47441 N47441 0 diode
R47442 N47441 N47442 10
D47442 N47442 0 diode
R47443 N47442 N47443 10
D47443 N47443 0 diode
R47444 N47443 N47444 10
D47444 N47444 0 diode
R47445 N47444 N47445 10
D47445 N47445 0 diode
R47446 N47445 N47446 10
D47446 N47446 0 diode
R47447 N47446 N47447 10
D47447 N47447 0 diode
R47448 N47447 N47448 10
D47448 N47448 0 diode
R47449 N47448 N47449 10
D47449 N47449 0 diode
R47450 N47449 N47450 10
D47450 N47450 0 diode
R47451 N47450 N47451 10
D47451 N47451 0 diode
R47452 N47451 N47452 10
D47452 N47452 0 diode
R47453 N47452 N47453 10
D47453 N47453 0 diode
R47454 N47453 N47454 10
D47454 N47454 0 diode
R47455 N47454 N47455 10
D47455 N47455 0 diode
R47456 N47455 N47456 10
D47456 N47456 0 diode
R47457 N47456 N47457 10
D47457 N47457 0 diode
R47458 N47457 N47458 10
D47458 N47458 0 diode
R47459 N47458 N47459 10
D47459 N47459 0 diode
R47460 N47459 N47460 10
D47460 N47460 0 diode
R47461 N47460 N47461 10
D47461 N47461 0 diode
R47462 N47461 N47462 10
D47462 N47462 0 diode
R47463 N47462 N47463 10
D47463 N47463 0 diode
R47464 N47463 N47464 10
D47464 N47464 0 diode
R47465 N47464 N47465 10
D47465 N47465 0 diode
R47466 N47465 N47466 10
D47466 N47466 0 diode
R47467 N47466 N47467 10
D47467 N47467 0 diode
R47468 N47467 N47468 10
D47468 N47468 0 diode
R47469 N47468 N47469 10
D47469 N47469 0 diode
R47470 N47469 N47470 10
D47470 N47470 0 diode
R47471 N47470 N47471 10
D47471 N47471 0 diode
R47472 N47471 N47472 10
D47472 N47472 0 diode
R47473 N47472 N47473 10
D47473 N47473 0 diode
R47474 N47473 N47474 10
D47474 N47474 0 diode
R47475 N47474 N47475 10
D47475 N47475 0 diode
R47476 N47475 N47476 10
D47476 N47476 0 diode
R47477 N47476 N47477 10
D47477 N47477 0 diode
R47478 N47477 N47478 10
D47478 N47478 0 diode
R47479 N47478 N47479 10
D47479 N47479 0 diode
R47480 N47479 N47480 10
D47480 N47480 0 diode
R47481 N47480 N47481 10
D47481 N47481 0 diode
R47482 N47481 N47482 10
D47482 N47482 0 diode
R47483 N47482 N47483 10
D47483 N47483 0 diode
R47484 N47483 N47484 10
D47484 N47484 0 diode
R47485 N47484 N47485 10
D47485 N47485 0 diode
R47486 N47485 N47486 10
D47486 N47486 0 diode
R47487 N47486 N47487 10
D47487 N47487 0 diode
R47488 N47487 N47488 10
D47488 N47488 0 diode
R47489 N47488 N47489 10
D47489 N47489 0 diode
R47490 N47489 N47490 10
D47490 N47490 0 diode
R47491 N47490 N47491 10
D47491 N47491 0 diode
R47492 N47491 N47492 10
D47492 N47492 0 diode
R47493 N47492 N47493 10
D47493 N47493 0 diode
R47494 N47493 N47494 10
D47494 N47494 0 diode
R47495 N47494 N47495 10
D47495 N47495 0 diode
R47496 N47495 N47496 10
D47496 N47496 0 diode
R47497 N47496 N47497 10
D47497 N47497 0 diode
R47498 N47497 N47498 10
D47498 N47498 0 diode
R47499 N47498 N47499 10
D47499 N47499 0 diode
R47500 N47499 N47500 10
D47500 N47500 0 diode
R47501 N47500 N47501 10
D47501 N47501 0 diode
R47502 N47501 N47502 10
D47502 N47502 0 diode
R47503 N47502 N47503 10
D47503 N47503 0 diode
R47504 N47503 N47504 10
D47504 N47504 0 diode
R47505 N47504 N47505 10
D47505 N47505 0 diode
R47506 N47505 N47506 10
D47506 N47506 0 diode
R47507 N47506 N47507 10
D47507 N47507 0 diode
R47508 N47507 N47508 10
D47508 N47508 0 diode
R47509 N47508 N47509 10
D47509 N47509 0 diode
R47510 N47509 N47510 10
D47510 N47510 0 diode
R47511 N47510 N47511 10
D47511 N47511 0 diode
R47512 N47511 N47512 10
D47512 N47512 0 diode
R47513 N47512 N47513 10
D47513 N47513 0 diode
R47514 N47513 N47514 10
D47514 N47514 0 diode
R47515 N47514 N47515 10
D47515 N47515 0 diode
R47516 N47515 N47516 10
D47516 N47516 0 diode
R47517 N47516 N47517 10
D47517 N47517 0 diode
R47518 N47517 N47518 10
D47518 N47518 0 diode
R47519 N47518 N47519 10
D47519 N47519 0 diode
R47520 N47519 N47520 10
D47520 N47520 0 diode
R47521 N47520 N47521 10
D47521 N47521 0 diode
R47522 N47521 N47522 10
D47522 N47522 0 diode
R47523 N47522 N47523 10
D47523 N47523 0 diode
R47524 N47523 N47524 10
D47524 N47524 0 diode
R47525 N47524 N47525 10
D47525 N47525 0 diode
R47526 N47525 N47526 10
D47526 N47526 0 diode
R47527 N47526 N47527 10
D47527 N47527 0 diode
R47528 N47527 N47528 10
D47528 N47528 0 diode
R47529 N47528 N47529 10
D47529 N47529 0 diode
R47530 N47529 N47530 10
D47530 N47530 0 diode
R47531 N47530 N47531 10
D47531 N47531 0 diode
R47532 N47531 N47532 10
D47532 N47532 0 diode
R47533 N47532 N47533 10
D47533 N47533 0 diode
R47534 N47533 N47534 10
D47534 N47534 0 diode
R47535 N47534 N47535 10
D47535 N47535 0 diode
R47536 N47535 N47536 10
D47536 N47536 0 diode
R47537 N47536 N47537 10
D47537 N47537 0 diode
R47538 N47537 N47538 10
D47538 N47538 0 diode
R47539 N47538 N47539 10
D47539 N47539 0 diode
R47540 N47539 N47540 10
D47540 N47540 0 diode
R47541 N47540 N47541 10
D47541 N47541 0 diode
R47542 N47541 N47542 10
D47542 N47542 0 diode
R47543 N47542 N47543 10
D47543 N47543 0 diode
R47544 N47543 N47544 10
D47544 N47544 0 diode
R47545 N47544 N47545 10
D47545 N47545 0 diode
R47546 N47545 N47546 10
D47546 N47546 0 diode
R47547 N47546 N47547 10
D47547 N47547 0 diode
R47548 N47547 N47548 10
D47548 N47548 0 diode
R47549 N47548 N47549 10
D47549 N47549 0 diode
R47550 N47549 N47550 10
D47550 N47550 0 diode
R47551 N47550 N47551 10
D47551 N47551 0 diode
R47552 N47551 N47552 10
D47552 N47552 0 diode
R47553 N47552 N47553 10
D47553 N47553 0 diode
R47554 N47553 N47554 10
D47554 N47554 0 diode
R47555 N47554 N47555 10
D47555 N47555 0 diode
R47556 N47555 N47556 10
D47556 N47556 0 diode
R47557 N47556 N47557 10
D47557 N47557 0 diode
R47558 N47557 N47558 10
D47558 N47558 0 diode
R47559 N47558 N47559 10
D47559 N47559 0 diode
R47560 N47559 N47560 10
D47560 N47560 0 diode
R47561 N47560 N47561 10
D47561 N47561 0 diode
R47562 N47561 N47562 10
D47562 N47562 0 diode
R47563 N47562 N47563 10
D47563 N47563 0 diode
R47564 N47563 N47564 10
D47564 N47564 0 diode
R47565 N47564 N47565 10
D47565 N47565 0 diode
R47566 N47565 N47566 10
D47566 N47566 0 diode
R47567 N47566 N47567 10
D47567 N47567 0 diode
R47568 N47567 N47568 10
D47568 N47568 0 diode
R47569 N47568 N47569 10
D47569 N47569 0 diode
R47570 N47569 N47570 10
D47570 N47570 0 diode
R47571 N47570 N47571 10
D47571 N47571 0 diode
R47572 N47571 N47572 10
D47572 N47572 0 diode
R47573 N47572 N47573 10
D47573 N47573 0 diode
R47574 N47573 N47574 10
D47574 N47574 0 diode
R47575 N47574 N47575 10
D47575 N47575 0 diode
R47576 N47575 N47576 10
D47576 N47576 0 diode
R47577 N47576 N47577 10
D47577 N47577 0 diode
R47578 N47577 N47578 10
D47578 N47578 0 diode
R47579 N47578 N47579 10
D47579 N47579 0 diode
R47580 N47579 N47580 10
D47580 N47580 0 diode
R47581 N47580 N47581 10
D47581 N47581 0 diode
R47582 N47581 N47582 10
D47582 N47582 0 diode
R47583 N47582 N47583 10
D47583 N47583 0 diode
R47584 N47583 N47584 10
D47584 N47584 0 diode
R47585 N47584 N47585 10
D47585 N47585 0 diode
R47586 N47585 N47586 10
D47586 N47586 0 diode
R47587 N47586 N47587 10
D47587 N47587 0 diode
R47588 N47587 N47588 10
D47588 N47588 0 diode
R47589 N47588 N47589 10
D47589 N47589 0 diode
R47590 N47589 N47590 10
D47590 N47590 0 diode
R47591 N47590 N47591 10
D47591 N47591 0 diode
R47592 N47591 N47592 10
D47592 N47592 0 diode
R47593 N47592 N47593 10
D47593 N47593 0 diode
R47594 N47593 N47594 10
D47594 N47594 0 diode
R47595 N47594 N47595 10
D47595 N47595 0 diode
R47596 N47595 N47596 10
D47596 N47596 0 diode
R47597 N47596 N47597 10
D47597 N47597 0 diode
R47598 N47597 N47598 10
D47598 N47598 0 diode
R47599 N47598 N47599 10
D47599 N47599 0 diode
R47600 N47599 N47600 10
D47600 N47600 0 diode
R47601 N47600 N47601 10
D47601 N47601 0 diode
R47602 N47601 N47602 10
D47602 N47602 0 diode
R47603 N47602 N47603 10
D47603 N47603 0 diode
R47604 N47603 N47604 10
D47604 N47604 0 diode
R47605 N47604 N47605 10
D47605 N47605 0 diode
R47606 N47605 N47606 10
D47606 N47606 0 diode
R47607 N47606 N47607 10
D47607 N47607 0 diode
R47608 N47607 N47608 10
D47608 N47608 0 diode
R47609 N47608 N47609 10
D47609 N47609 0 diode
R47610 N47609 N47610 10
D47610 N47610 0 diode
R47611 N47610 N47611 10
D47611 N47611 0 diode
R47612 N47611 N47612 10
D47612 N47612 0 diode
R47613 N47612 N47613 10
D47613 N47613 0 diode
R47614 N47613 N47614 10
D47614 N47614 0 diode
R47615 N47614 N47615 10
D47615 N47615 0 diode
R47616 N47615 N47616 10
D47616 N47616 0 diode
R47617 N47616 N47617 10
D47617 N47617 0 diode
R47618 N47617 N47618 10
D47618 N47618 0 diode
R47619 N47618 N47619 10
D47619 N47619 0 diode
R47620 N47619 N47620 10
D47620 N47620 0 diode
R47621 N47620 N47621 10
D47621 N47621 0 diode
R47622 N47621 N47622 10
D47622 N47622 0 diode
R47623 N47622 N47623 10
D47623 N47623 0 diode
R47624 N47623 N47624 10
D47624 N47624 0 diode
R47625 N47624 N47625 10
D47625 N47625 0 diode
R47626 N47625 N47626 10
D47626 N47626 0 diode
R47627 N47626 N47627 10
D47627 N47627 0 diode
R47628 N47627 N47628 10
D47628 N47628 0 diode
R47629 N47628 N47629 10
D47629 N47629 0 diode
R47630 N47629 N47630 10
D47630 N47630 0 diode
R47631 N47630 N47631 10
D47631 N47631 0 diode
R47632 N47631 N47632 10
D47632 N47632 0 diode
R47633 N47632 N47633 10
D47633 N47633 0 diode
R47634 N47633 N47634 10
D47634 N47634 0 diode
R47635 N47634 N47635 10
D47635 N47635 0 diode
R47636 N47635 N47636 10
D47636 N47636 0 diode
R47637 N47636 N47637 10
D47637 N47637 0 diode
R47638 N47637 N47638 10
D47638 N47638 0 diode
R47639 N47638 N47639 10
D47639 N47639 0 diode
R47640 N47639 N47640 10
D47640 N47640 0 diode
R47641 N47640 N47641 10
D47641 N47641 0 diode
R47642 N47641 N47642 10
D47642 N47642 0 diode
R47643 N47642 N47643 10
D47643 N47643 0 diode
R47644 N47643 N47644 10
D47644 N47644 0 diode
R47645 N47644 N47645 10
D47645 N47645 0 diode
R47646 N47645 N47646 10
D47646 N47646 0 diode
R47647 N47646 N47647 10
D47647 N47647 0 diode
R47648 N47647 N47648 10
D47648 N47648 0 diode
R47649 N47648 N47649 10
D47649 N47649 0 diode
R47650 N47649 N47650 10
D47650 N47650 0 diode
R47651 N47650 N47651 10
D47651 N47651 0 diode
R47652 N47651 N47652 10
D47652 N47652 0 diode
R47653 N47652 N47653 10
D47653 N47653 0 diode
R47654 N47653 N47654 10
D47654 N47654 0 diode
R47655 N47654 N47655 10
D47655 N47655 0 diode
R47656 N47655 N47656 10
D47656 N47656 0 diode
R47657 N47656 N47657 10
D47657 N47657 0 diode
R47658 N47657 N47658 10
D47658 N47658 0 diode
R47659 N47658 N47659 10
D47659 N47659 0 diode
R47660 N47659 N47660 10
D47660 N47660 0 diode
R47661 N47660 N47661 10
D47661 N47661 0 diode
R47662 N47661 N47662 10
D47662 N47662 0 diode
R47663 N47662 N47663 10
D47663 N47663 0 diode
R47664 N47663 N47664 10
D47664 N47664 0 diode
R47665 N47664 N47665 10
D47665 N47665 0 diode
R47666 N47665 N47666 10
D47666 N47666 0 diode
R47667 N47666 N47667 10
D47667 N47667 0 diode
R47668 N47667 N47668 10
D47668 N47668 0 diode
R47669 N47668 N47669 10
D47669 N47669 0 diode
R47670 N47669 N47670 10
D47670 N47670 0 diode
R47671 N47670 N47671 10
D47671 N47671 0 diode
R47672 N47671 N47672 10
D47672 N47672 0 diode
R47673 N47672 N47673 10
D47673 N47673 0 diode
R47674 N47673 N47674 10
D47674 N47674 0 diode
R47675 N47674 N47675 10
D47675 N47675 0 diode
R47676 N47675 N47676 10
D47676 N47676 0 diode
R47677 N47676 N47677 10
D47677 N47677 0 diode
R47678 N47677 N47678 10
D47678 N47678 0 diode
R47679 N47678 N47679 10
D47679 N47679 0 diode
R47680 N47679 N47680 10
D47680 N47680 0 diode
R47681 N47680 N47681 10
D47681 N47681 0 diode
R47682 N47681 N47682 10
D47682 N47682 0 diode
R47683 N47682 N47683 10
D47683 N47683 0 diode
R47684 N47683 N47684 10
D47684 N47684 0 diode
R47685 N47684 N47685 10
D47685 N47685 0 diode
R47686 N47685 N47686 10
D47686 N47686 0 diode
R47687 N47686 N47687 10
D47687 N47687 0 diode
R47688 N47687 N47688 10
D47688 N47688 0 diode
R47689 N47688 N47689 10
D47689 N47689 0 diode
R47690 N47689 N47690 10
D47690 N47690 0 diode
R47691 N47690 N47691 10
D47691 N47691 0 diode
R47692 N47691 N47692 10
D47692 N47692 0 diode
R47693 N47692 N47693 10
D47693 N47693 0 diode
R47694 N47693 N47694 10
D47694 N47694 0 diode
R47695 N47694 N47695 10
D47695 N47695 0 diode
R47696 N47695 N47696 10
D47696 N47696 0 diode
R47697 N47696 N47697 10
D47697 N47697 0 diode
R47698 N47697 N47698 10
D47698 N47698 0 diode
R47699 N47698 N47699 10
D47699 N47699 0 diode
R47700 N47699 N47700 10
D47700 N47700 0 diode
R47701 N47700 N47701 10
D47701 N47701 0 diode
R47702 N47701 N47702 10
D47702 N47702 0 diode
R47703 N47702 N47703 10
D47703 N47703 0 diode
R47704 N47703 N47704 10
D47704 N47704 0 diode
R47705 N47704 N47705 10
D47705 N47705 0 diode
R47706 N47705 N47706 10
D47706 N47706 0 diode
R47707 N47706 N47707 10
D47707 N47707 0 diode
R47708 N47707 N47708 10
D47708 N47708 0 diode
R47709 N47708 N47709 10
D47709 N47709 0 diode
R47710 N47709 N47710 10
D47710 N47710 0 diode
R47711 N47710 N47711 10
D47711 N47711 0 diode
R47712 N47711 N47712 10
D47712 N47712 0 diode
R47713 N47712 N47713 10
D47713 N47713 0 diode
R47714 N47713 N47714 10
D47714 N47714 0 diode
R47715 N47714 N47715 10
D47715 N47715 0 diode
R47716 N47715 N47716 10
D47716 N47716 0 diode
R47717 N47716 N47717 10
D47717 N47717 0 diode
R47718 N47717 N47718 10
D47718 N47718 0 diode
R47719 N47718 N47719 10
D47719 N47719 0 diode
R47720 N47719 N47720 10
D47720 N47720 0 diode
R47721 N47720 N47721 10
D47721 N47721 0 diode
R47722 N47721 N47722 10
D47722 N47722 0 diode
R47723 N47722 N47723 10
D47723 N47723 0 diode
R47724 N47723 N47724 10
D47724 N47724 0 diode
R47725 N47724 N47725 10
D47725 N47725 0 diode
R47726 N47725 N47726 10
D47726 N47726 0 diode
R47727 N47726 N47727 10
D47727 N47727 0 diode
R47728 N47727 N47728 10
D47728 N47728 0 diode
R47729 N47728 N47729 10
D47729 N47729 0 diode
R47730 N47729 N47730 10
D47730 N47730 0 diode
R47731 N47730 N47731 10
D47731 N47731 0 diode
R47732 N47731 N47732 10
D47732 N47732 0 diode
R47733 N47732 N47733 10
D47733 N47733 0 diode
R47734 N47733 N47734 10
D47734 N47734 0 diode
R47735 N47734 N47735 10
D47735 N47735 0 diode
R47736 N47735 N47736 10
D47736 N47736 0 diode
R47737 N47736 N47737 10
D47737 N47737 0 diode
R47738 N47737 N47738 10
D47738 N47738 0 diode
R47739 N47738 N47739 10
D47739 N47739 0 diode
R47740 N47739 N47740 10
D47740 N47740 0 diode
R47741 N47740 N47741 10
D47741 N47741 0 diode
R47742 N47741 N47742 10
D47742 N47742 0 diode
R47743 N47742 N47743 10
D47743 N47743 0 diode
R47744 N47743 N47744 10
D47744 N47744 0 diode
R47745 N47744 N47745 10
D47745 N47745 0 diode
R47746 N47745 N47746 10
D47746 N47746 0 diode
R47747 N47746 N47747 10
D47747 N47747 0 diode
R47748 N47747 N47748 10
D47748 N47748 0 diode
R47749 N47748 N47749 10
D47749 N47749 0 diode
R47750 N47749 N47750 10
D47750 N47750 0 diode
R47751 N47750 N47751 10
D47751 N47751 0 diode
R47752 N47751 N47752 10
D47752 N47752 0 diode
R47753 N47752 N47753 10
D47753 N47753 0 diode
R47754 N47753 N47754 10
D47754 N47754 0 diode
R47755 N47754 N47755 10
D47755 N47755 0 diode
R47756 N47755 N47756 10
D47756 N47756 0 diode
R47757 N47756 N47757 10
D47757 N47757 0 diode
R47758 N47757 N47758 10
D47758 N47758 0 diode
R47759 N47758 N47759 10
D47759 N47759 0 diode
R47760 N47759 N47760 10
D47760 N47760 0 diode
R47761 N47760 N47761 10
D47761 N47761 0 diode
R47762 N47761 N47762 10
D47762 N47762 0 diode
R47763 N47762 N47763 10
D47763 N47763 0 diode
R47764 N47763 N47764 10
D47764 N47764 0 diode
R47765 N47764 N47765 10
D47765 N47765 0 diode
R47766 N47765 N47766 10
D47766 N47766 0 diode
R47767 N47766 N47767 10
D47767 N47767 0 diode
R47768 N47767 N47768 10
D47768 N47768 0 diode
R47769 N47768 N47769 10
D47769 N47769 0 diode
R47770 N47769 N47770 10
D47770 N47770 0 diode
R47771 N47770 N47771 10
D47771 N47771 0 diode
R47772 N47771 N47772 10
D47772 N47772 0 diode
R47773 N47772 N47773 10
D47773 N47773 0 diode
R47774 N47773 N47774 10
D47774 N47774 0 diode
R47775 N47774 N47775 10
D47775 N47775 0 diode
R47776 N47775 N47776 10
D47776 N47776 0 diode
R47777 N47776 N47777 10
D47777 N47777 0 diode
R47778 N47777 N47778 10
D47778 N47778 0 diode
R47779 N47778 N47779 10
D47779 N47779 0 diode
R47780 N47779 N47780 10
D47780 N47780 0 diode
R47781 N47780 N47781 10
D47781 N47781 0 diode
R47782 N47781 N47782 10
D47782 N47782 0 diode
R47783 N47782 N47783 10
D47783 N47783 0 diode
R47784 N47783 N47784 10
D47784 N47784 0 diode
R47785 N47784 N47785 10
D47785 N47785 0 diode
R47786 N47785 N47786 10
D47786 N47786 0 diode
R47787 N47786 N47787 10
D47787 N47787 0 diode
R47788 N47787 N47788 10
D47788 N47788 0 diode
R47789 N47788 N47789 10
D47789 N47789 0 diode
R47790 N47789 N47790 10
D47790 N47790 0 diode
R47791 N47790 N47791 10
D47791 N47791 0 diode
R47792 N47791 N47792 10
D47792 N47792 0 diode
R47793 N47792 N47793 10
D47793 N47793 0 diode
R47794 N47793 N47794 10
D47794 N47794 0 diode
R47795 N47794 N47795 10
D47795 N47795 0 diode
R47796 N47795 N47796 10
D47796 N47796 0 diode
R47797 N47796 N47797 10
D47797 N47797 0 diode
R47798 N47797 N47798 10
D47798 N47798 0 diode
R47799 N47798 N47799 10
D47799 N47799 0 diode
R47800 N47799 N47800 10
D47800 N47800 0 diode
R47801 N47800 N47801 10
D47801 N47801 0 diode
R47802 N47801 N47802 10
D47802 N47802 0 diode
R47803 N47802 N47803 10
D47803 N47803 0 diode
R47804 N47803 N47804 10
D47804 N47804 0 diode
R47805 N47804 N47805 10
D47805 N47805 0 diode
R47806 N47805 N47806 10
D47806 N47806 0 diode
R47807 N47806 N47807 10
D47807 N47807 0 diode
R47808 N47807 N47808 10
D47808 N47808 0 diode
R47809 N47808 N47809 10
D47809 N47809 0 diode
R47810 N47809 N47810 10
D47810 N47810 0 diode
R47811 N47810 N47811 10
D47811 N47811 0 diode
R47812 N47811 N47812 10
D47812 N47812 0 diode
R47813 N47812 N47813 10
D47813 N47813 0 diode
R47814 N47813 N47814 10
D47814 N47814 0 diode
R47815 N47814 N47815 10
D47815 N47815 0 diode
R47816 N47815 N47816 10
D47816 N47816 0 diode
R47817 N47816 N47817 10
D47817 N47817 0 diode
R47818 N47817 N47818 10
D47818 N47818 0 diode
R47819 N47818 N47819 10
D47819 N47819 0 diode
R47820 N47819 N47820 10
D47820 N47820 0 diode
R47821 N47820 N47821 10
D47821 N47821 0 diode
R47822 N47821 N47822 10
D47822 N47822 0 diode
R47823 N47822 N47823 10
D47823 N47823 0 diode
R47824 N47823 N47824 10
D47824 N47824 0 diode
R47825 N47824 N47825 10
D47825 N47825 0 diode
R47826 N47825 N47826 10
D47826 N47826 0 diode
R47827 N47826 N47827 10
D47827 N47827 0 diode
R47828 N47827 N47828 10
D47828 N47828 0 diode
R47829 N47828 N47829 10
D47829 N47829 0 diode
R47830 N47829 N47830 10
D47830 N47830 0 diode
R47831 N47830 N47831 10
D47831 N47831 0 diode
R47832 N47831 N47832 10
D47832 N47832 0 diode
R47833 N47832 N47833 10
D47833 N47833 0 diode
R47834 N47833 N47834 10
D47834 N47834 0 diode
R47835 N47834 N47835 10
D47835 N47835 0 diode
R47836 N47835 N47836 10
D47836 N47836 0 diode
R47837 N47836 N47837 10
D47837 N47837 0 diode
R47838 N47837 N47838 10
D47838 N47838 0 diode
R47839 N47838 N47839 10
D47839 N47839 0 diode
R47840 N47839 N47840 10
D47840 N47840 0 diode
R47841 N47840 N47841 10
D47841 N47841 0 diode
R47842 N47841 N47842 10
D47842 N47842 0 diode
R47843 N47842 N47843 10
D47843 N47843 0 diode
R47844 N47843 N47844 10
D47844 N47844 0 diode
R47845 N47844 N47845 10
D47845 N47845 0 diode
R47846 N47845 N47846 10
D47846 N47846 0 diode
R47847 N47846 N47847 10
D47847 N47847 0 diode
R47848 N47847 N47848 10
D47848 N47848 0 diode
R47849 N47848 N47849 10
D47849 N47849 0 diode
R47850 N47849 N47850 10
D47850 N47850 0 diode
R47851 N47850 N47851 10
D47851 N47851 0 diode
R47852 N47851 N47852 10
D47852 N47852 0 diode
R47853 N47852 N47853 10
D47853 N47853 0 diode
R47854 N47853 N47854 10
D47854 N47854 0 diode
R47855 N47854 N47855 10
D47855 N47855 0 diode
R47856 N47855 N47856 10
D47856 N47856 0 diode
R47857 N47856 N47857 10
D47857 N47857 0 diode
R47858 N47857 N47858 10
D47858 N47858 0 diode
R47859 N47858 N47859 10
D47859 N47859 0 diode
R47860 N47859 N47860 10
D47860 N47860 0 diode
R47861 N47860 N47861 10
D47861 N47861 0 diode
R47862 N47861 N47862 10
D47862 N47862 0 diode
R47863 N47862 N47863 10
D47863 N47863 0 diode
R47864 N47863 N47864 10
D47864 N47864 0 diode
R47865 N47864 N47865 10
D47865 N47865 0 diode
R47866 N47865 N47866 10
D47866 N47866 0 diode
R47867 N47866 N47867 10
D47867 N47867 0 diode
R47868 N47867 N47868 10
D47868 N47868 0 diode
R47869 N47868 N47869 10
D47869 N47869 0 diode
R47870 N47869 N47870 10
D47870 N47870 0 diode
R47871 N47870 N47871 10
D47871 N47871 0 diode
R47872 N47871 N47872 10
D47872 N47872 0 diode
R47873 N47872 N47873 10
D47873 N47873 0 diode
R47874 N47873 N47874 10
D47874 N47874 0 diode
R47875 N47874 N47875 10
D47875 N47875 0 diode
R47876 N47875 N47876 10
D47876 N47876 0 diode
R47877 N47876 N47877 10
D47877 N47877 0 diode
R47878 N47877 N47878 10
D47878 N47878 0 diode
R47879 N47878 N47879 10
D47879 N47879 0 diode
R47880 N47879 N47880 10
D47880 N47880 0 diode
R47881 N47880 N47881 10
D47881 N47881 0 diode
R47882 N47881 N47882 10
D47882 N47882 0 diode
R47883 N47882 N47883 10
D47883 N47883 0 diode
R47884 N47883 N47884 10
D47884 N47884 0 diode
R47885 N47884 N47885 10
D47885 N47885 0 diode
R47886 N47885 N47886 10
D47886 N47886 0 diode
R47887 N47886 N47887 10
D47887 N47887 0 diode
R47888 N47887 N47888 10
D47888 N47888 0 diode
R47889 N47888 N47889 10
D47889 N47889 0 diode
R47890 N47889 N47890 10
D47890 N47890 0 diode
R47891 N47890 N47891 10
D47891 N47891 0 diode
R47892 N47891 N47892 10
D47892 N47892 0 diode
R47893 N47892 N47893 10
D47893 N47893 0 diode
R47894 N47893 N47894 10
D47894 N47894 0 diode
R47895 N47894 N47895 10
D47895 N47895 0 diode
R47896 N47895 N47896 10
D47896 N47896 0 diode
R47897 N47896 N47897 10
D47897 N47897 0 diode
R47898 N47897 N47898 10
D47898 N47898 0 diode
R47899 N47898 N47899 10
D47899 N47899 0 diode
R47900 N47899 N47900 10
D47900 N47900 0 diode
R47901 N47900 N47901 10
D47901 N47901 0 diode
R47902 N47901 N47902 10
D47902 N47902 0 diode
R47903 N47902 N47903 10
D47903 N47903 0 diode
R47904 N47903 N47904 10
D47904 N47904 0 diode
R47905 N47904 N47905 10
D47905 N47905 0 diode
R47906 N47905 N47906 10
D47906 N47906 0 diode
R47907 N47906 N47907 10
D47907 N47907 0 diode
R47908 N47907 N47908 10
D47908 N47908 0 diode
R47909 N47908 N47909 10
D47909 N47909 0 diode
R47910 N47909 N47910 10
D47910 N47910 0 diode
R47911 N47910 N47911 10
D47911 N47911 0 diode
R47912 N47911 N47912 10
D47912 N47912 0 diode
R47913 N47912 N47913 10
D47913 N47913 0 diode
R47914 N47913 N47914 10
D47914 N47914 0 diode
R47915 N47914 N47915 10
D47915 N47915 0 diode
R47916 N47915 N47916 10
D47916 N47916 0 diode
R47917 N47916 N47917 10
D47917 N47917 0 diode
R47918 N47917 N47918 10
D47918 N47918 0 diode
R47919 N47918 N47919 10
D47919 N47919 0 diode
R47920 N47919 N47920 10
D47920 N47920 0 diode
R47921 N47920 N47921 10
D47921 N47921 0 diode
R47922 N47921 N47922 10
D47922 N47922 0 diode
R47923 N47922 N47923 10
D47923 N47923 0 diode
R47924 N47923 N47924 10
D47924 N47924 0 diode
R47925 N47924 N47925 10
D47925 N47925 0 diode
R47926 N47925 N47926 10
D47926 N47926 0 diode
R47927 N47926 N47927 10
D47927 N47927 0 diode
R47928 N47927 N47928 10
D47928 N47928 0 diode
R47929 N47928 N47929 10
D47929 N47929 0 diode
R47930 N47929 N47930 10
D47930 N47930 0 diode
R47931 N47930 N47931 10
D47931 N47931 0 diode
R47932 N47931 N47932 10
D47932 N47932 0 diode
R47933 N47932 N47933 10
D47933 N47933 0 diode
R47934 N47933 N47934 10
D47934 N47934 0 diode
R47935 N47934 N47935 10
D47935 N47935 0 diode
R47936 N47935 N47936 10
D47936 N47936 0 diode
R47937 N47936 N47937 10
D47937 N47937 0 diode
R47938 N47937 N47938 10
D47938 N47938 0 diode
R47939 N47938 N47939 10
D47939 N47939 0 diode
R47940 N47939 N47940 10
D47940 N47940 0 diode
R47941 N47940 N47941 10
D47941 N47941 0 diode
R47942 N47941 N47942 10
D47942 N47942 0 diode
R47943 N47942 N47943 10
D47943 N47943 0 diode
R47944 N47943 N47944 10
D47944 N47944 0 diode
R47945 N47944 N47945 10
D47945 N47945 0 diode
R47946 N47945 N47946 10
D47946 N47946 0 diode
R47947 N47946 N47947 10
D47947 N47947 0 diode
R47948 N47947 N47948 10
D47948 N47948 0 diode
R47949 N47948 N47949 10
D47949 N47949 0 diode
R47950 N47949 N47950 10
D47950 N47950 0 diode
R47951 N47950 N47951 10
D47951 N47951 0 diode
R47952 N47951 N47952 10
D47952 N47952 0 diode
R47953 N47952 N47953 10
D47953 N47953 0 diode
R47954 N47953 N47954 10
D47954 N47954 0 diode
R47955 N47954 N47955 10
D47955 N47955 0 diode
R47956 N47955 N47956 10
D47956 N47956 0 diode
R47957 N47956 N47957 10
D47957 N47957 0 diode
R47958 N47957 N47958 10
D47958 N47958 0 diode
R47959 N47958 N47959 10
D47959 N47959 0 diode
R47960 N47959 N47960 10
D47960 N47960 0 diode
R47961 N47960 N47961 10
D47961 N47961 0 diode
R47962 N47961 N47962 10
D47962 N47962 0 diode
R47963 N47962 N47963 10
D47963 N47963 0 diode
R47964 N47963 N47964 10
D47964 N47964 0 diode
R47965 N47964 N47965 10
D47965 N47965 0 diode
R47966 N47965 N47966 10
D47966 N47966 0 diode
R47967 N47966 N47967 10
D47967 N47967 0 diode
R47968 N47967 N47968 10
D47968 N47968 0 diode
R47969 N47968 N47969 10
D47969 N47969 0 diode
R47970 N47969 N47970 10
D47970 N47970 0 diode
R47971 N47970 N47971 10
D47971 N47971 0 diode
R47972 N47971 N47972 10
D47972 N47972 0 diode
R47973 N47972 N47973 10
D47973 N47973 0 diode
R47974 N47973 N47974 10
D47974 N47974 0 diode
R47975 N47974 N47975 10
D47975 N47975 0 diode
R47976 N47975 N47976 10
D47976 N47976 0 diode
R47977 N47976 N47977 10
D47977 N47977 0 diode
R47978 N47977 N47978 10
D47978 N47978 0 diode
R47979 N47978 N47979 10
D47979 N47979 0 diode
R47980 N47979 N47980 10
D47980 N47980 0 diode
R47981 N47980 N47981 10
D47981 N47981 0 diode
R47982 N47981 N47982 10
D47982 N47982 0 diode
R47983 N47982 N47983 10
D47983 N47983 0 diode
R47984 N47983 N47984 10
D47984 N47984 0 diode
R47985 N47984 N47985 10
D47985 N47985 0 diode
R47986 N47985 N47986 10
D47986 N47986 0 diode
R47987 N47986 N47987 10
D47987 N47987 0 diode
R47988 N47987 N47988 10
D47988 N47988 0 diode
R47989 N47988 N47989 10
D47989 N47989 0 diode
R47990 N47989 N47990 10
D47990 N47990 0 diode
R47991 N47990 N47991 10
D47991 N47991 0 diode
R47992 N47991 N47992 10
D47992 N47992 0 diode
R47993 N47992 N47993 10
D47993 N47993 0 diode
R47994 N47993 N47994 10
D47994 N47994 0 diode
R47995 N47994 N47995 10
D47995 N47995 0 diode
R47996 N47995 N47996 10
D47996 N47996 0 diode
R47997 N47996 N47997 10
D47997 N47997 0 diode
R47998 N47997 N47998 10
D47998 N47998 0 diode
R47999 N47998 N47999 10
D47999 N47999 0 diode
R48000 N47999 N48000 10
D48000 N48000 0 diode
R48001 N48000 N48001 10
D48001 N48001 0 diode
R48002 N48001 N48002 10
D48002 N48002 0 diode
R48003 N48002 N48003 10
D48003 N48003 0 diode
R48004 N48003 N48004 10
D48004 N48004 0 diode
R48005 N48004 N48005 10
D48005 N48005 0 diode
R48006 N48005 N48006 10
D48006 N48006 0 diode
R48007 N48006 N48007 10
D48007 N48007 0 diode
R48008 N48007 N48008 10
D48008 N48008 0 diode
R48009 N48008 N48009 10
D48009 N48009 0 diode
R48010 N48009 N48010 10
D48010 N48010 0 diode
R48011 N48010 N48011 10
D48011 N48011 0 diode
R48012 N48011 N48012 10
D48012 N48012 0 diode
R48013 N48012 N48013 10
D48013 N48013 0 diode
R48014 N48013 N48014 10
D48014 N48014 0 diode
R48015 N48014 N48015 10
D48015 N48015 0 diode
R48016 N48015 N48016 10
D48016 N48016 0 diode
R48017 N48016 N48017 10
D48017 N48017 0 diode
R48018 N48017 N48018 10
D48018 N48018 0 diode
R48019 N48018 N48019 10
D48019 N48019 0 diode
R48020 N48019 N48020 10
D48020 N48020 0 diode
R48021 N48020 N48021 10
D48021 N48021 0 diode
R48022 N48021 N48022 10
D48022 N48022 0 diode
R48023 N48022 N48023 10
D48023 N48023 0 diode
R48024 N48023 N48024 10
D48024 N48024 0 diode
R48025 N48024 N48025 10
D48025 N48025 0 diode
R48026 N48025 N48026 10
D48026 N48026 0 diode
R48027 N48026 N48027 10
D48027 N48027 0 diode
R48028 N48027 N48028 10
D48028 N48028 0 diode
R48029 N48028 N48029 10
D48029 N48029 0 diode
R48030 N48029 N48030 10
D48030 N48030 0 diode
R48031 N48030 N48031 10
D48031 N48031 0 diode
R48032 N48031 N48032 10
D48032 N48032 0 diode
R48033 N48032 N48033 10
D48033 N48033 0 diode
R48034 N48033 N48034 10
D48034 N48034 0 diode
R48035 N48034 N48035 10
D48035 N48035 0 diode
R48036 N48035 N48036 10
D48036 N48036 0 diode
R48037 N48036 N48037 10
D48037 N48037 0 diode
R48038 N48037 N48038 10
D48038 N48038 0 diode
R48039 N48038 N48039 10
D48039 N48039 0 diode
R48040 N48039 N48040 10
D48040 N48040 0 diode
R48041 N48040 N48041 10
D48041 N48041 0 diode
R48042 N48041 N48042 10
D48042 N48042 0 diode
R48043 N48042 N48043 10
D48043 N48043 0 diode
R48044 N48043 N48044 10
D48044 N48044 0 diode
R48045 N48044 N48045 10
D48045 N48045 0 diode
R48046 N48045 N48046 10
D48046 N48046 0 diode
R48047 N48046 N48047 10
D48047 N48047 0 diode
R48048 N48047 N48048 10
D48048 N48048 0 diode
R48049 N48048 N48049 10
D48049 N48049 0 diode
R48050 N48049 N48050 10
D48050 N48050 0 diode
R48051 N48050 N48051 10
D48051 N48051 0 diode
R48052 N48051 N48052 10
D48052 N48052 0 diode
R48053 N48052 N48053 10
D48053 N48053 0 diode
R48054 N48053 N48054 10
D48054 N48054 0 diode
R48055 N48054 N48055 10
D48055 N48055 0 diode
R48056 N48055 N48056 10
D48056 N48056 0 diode
R48057 N48056 N48057 10
D48057 N48057 0 diode
R48058 N48057 N48058 10
D48058 N48058 0 diode
R48059 N48058 N48059 10
D48059 N48059 0 diode
R48060 N48059 N48060 10
D48060 N48060 0 diode
R48061 N48060 N48061 10
D48061 N48061 0 diode
R48062 N48061 N48062 10
D48062 N48062 0 diode
R48063 N48062 N48063 10
D48063 N48063 0 diode
R48064 N48063 N48064 10
D48064 N48064 0 diode
R48065 N48064 N48065 10
D48065 N48065 0 diode
R48066 N48065 N48066 10
D48066 N48066 0 diode
R48067 N48066 N48067 10
D48067 N48067 0 diode
R48068 N48067 N48068 10
D48068 N48068 0 diode
R48069 N48068 N48069 10
D48069 N48069 0 diode
R48070 N48069 N48070 10
D48070 N48070 0 diode
R48071 N48070 N48071 10
D48071 N48071 0 diode
R48072 N48071 N48072 10
D48072 N48072 0 diode
R48073 N48072 N48073 10
D48073 N48073 0 diode
R48074 N48073 N48074 10
D48074 N48074 0 diode
R48075 N48074 N48075 10
D48075 N48075 0 diode
R48076 N48075 N48076 10
D48076 N48076 0 diode
R48077 N48076 N48077 10
D48077 N48077 0 diode
R48078 N48077 N48078 10
D48078 N48078 0 diode
R48079 N48078 N48079 10
D48079 N48079 0 diode
R48080 N48079 N48080 10
D48080 N48080 0 diode
R48081 N48080 N48081 10
D48081 N48081 0 diode
R48082 N48081 N48082 10
D48082 N48082 0 diode
R48083 N48082 N48083 10
D48083 N48083 0 diode
R48084 N48083 N48084 10
D48084 N48084 0 diode
R48085 N48084 N48085 10
D48085 N48085 0 diode
R48086 N48085 N48086 10
D48086 N48086 0 diode
R48087 N48086 N48087 10
D48087 N48087 0 diode
R48088 N48087 N48088 10
D48088 N48088 0 diode
R48089 N48088 N48089 10
D48089 N48089 0 diode
R48090 N48089 N48090 10
D48090 N48090 0 diode
R48091 N48090 N48091 10
D48091 N48091 0 diode
R48092 N48091 N48092 10
D48092 N48092 0 diode
R48093 N48092 N48093 10
D48093 N48093 0 diode
R48094 N48093 N48094 10
D48094 N48094 0 diode
R48095 N48094 N48095 10
D48095 N48095 0 diode
R48096 N48095 N48096 10
D48096 N48096 0 diode
R48097 N48096 N48097 10
D48097 N48097 0 diode
R48098 N48097 N48098 10
D48098 N48098 0 diode
R48099 N48098 N48099 10
D48099 N48099 0 diode
R48100 N48099 N48100 10
D48100 N48100 0 diode
R48101 N48100 N48101 10
D48101 N48101 0 diode
R48102 N48101 N48102 10
D48102 N48102 0 diode
R48103 N48102 N48103 10
D48103 N48103 0 diode
R48104 N48103 N48104 10
D48104 N48104 0 diode
R48105 N48104 N48105 10
D48105 N48105 0 diode
R48106 N48105 N48106 10
D48106 N48106 0 diode
R48107 N48106 N48107 10
D48107 N48107 0 diode
R48108 N48107 N48108 10
D48108 N48108 0 diode
R48109 N48108 N48109 10
D48109 N48109 0 diode
R48110 N48109 N48110 10
D48110 N48110 0 diode
R48111 N48110 N48111 10
D48111 N48111 0 diode
R48112 N48111 N48112 10
D48112 N48112 0 diode
R48113 N48112 N48113 10
D48113 N48113 0 diode
R48114 N48113 N48114 10
D48114 N48114 0 diode
R48115 N48114 N48115 10
D48115 N48115 0 diode
R48116 N48115 N48116 10
D48116 N48116 0 diode
R48117 N48116 N48117 10
D48117 N48117 0 diode
R48118 N48117 N48118 10
D48118 N48118 0 diode
R48119 N48118 N48119 10
D48119 N48119 0 diode
R48120 N48119 N48120 10
D48120 N48120 0 diode
R48121 N48120 N48121 10
D48121 N48121 0 diode
R48122 N48121 N48122 10
D48122 N48122 0 diode
R48123 N48122 N48123 10
D48123 N48123 0 diode
R48124 N48123 N48124 10
D48124 N48124 0 diode
R48125 N48124 N48125 10
D48125 N48125 0 diode
R48126 N48125 N48126 10
D48126 N48126 0 diode
R48127 N48126 N48127 10
D48127 N48127 0 diode
R48128 N48127 N48128 10
D48128 N48128 0 diode
R48129 N48128 N48129 10
D48129 N48129 0 diode
R48130 N48129 N48130 10
D48130 N48130 0 diode
R48131 N48130 N48131 10
D48131 N48131 0 diode
R48132 N48131 N48132 10
D48132 N48132 0 diode
R48133 N48132 N48133 10
D48133 N48133 0 diode
R48134 N48133 N48134 10
D48134 N48134 0 diode
R48135 N48134 N48135 10
D48135 N48135 0 diode
R48136 N48135 N48136 10
D48136 N48136 0 diode
R48137 N48136 N48137 10
D48137 N48137 0 diode
R48138 N48137 N48138 10
D48138 N48138 0 diode
R48139 N48138 N48139 10
D48139 N48139 0 diode
R48140 N48139 N48140 10
D48140 N48140 0 diode
R48141 N48140 N48141 10
D48141 N48141 0 diode
R48142 N48141 N48142 10
D48142 N48142 0 diode
R48143 N48142 N48143 10
D48143 N48143 0 diode
R48144 N48143 N48144 10
D48144 N48144 0 diode
R48145 N48144 N48145 10
D48145 N48145 0 diode
R48146 N48145 N48146 10
D48146 N48146 0 diode
R48147 N48146 N48147 10
D48147 N48147 0 diode
R48148 N48147 N48148 10
D48148 N48148 0 diode
R48149 N48148 N48149 10
D48149 N48149 0 diode
R48150 N48149 N48150 10
D48150 N48150 0 diode
R48151 N48150 N48151 10
D48151 N48151 0 diode
R48152 N48151 N48152 10
D48152 N48152 0 diode
R48153 N48152 N48153 10
D48153 N48153 0 diode
R48154 N48153 N48154 10
D48154 N48154 0 diode
R48155 N48154 N48155 10
D48155 N48155 0 diode
R48156 N48155 N48156 10
D48156 N48156 0 diode
R48157 N48156 N48157 10
D48157 N48157 0 diode
R48158 N48157 N48158 10
D48158 N48158 0 diode
R48159 N48158 N48159 10
D48159 N48159 0 diode
R48160 N48159 N48160 10
D48160 N48160 0 diode
R48161 N48160 N48161 10
D48161 N48161 0 diode
R48162 N48161 N48162 10
D48162 N48162 0 diode
R48163 N48162 N48163 10
D48163 N48163 0 diode
R48164 N48163 N48164 10
D48164 N48164 0 diode
R48165 N48164 N48165 10
D48165 N48165 0 diode
R48166 N48165 N48166 10
D48166 N48166 0 diode
R48167 N48166 N48167 10
D48167 N48167 0 diode
R48168 N48167 N48168 10
D48168 N48168 0 diode
R48169 N48168 N48169 10
D48169 N48169 0 diode
R48170 N48169 N48170 10
D48170 N48170 0 diode
R48171 N48170 N48171 10
D48171 N48171 0 diode
R48172 N48171 N48172 10
D48172 N48172 0 diode
R48173 N48172 N48173 10
D48173 N48173 0 diode
R48174 N48173 N48174 10
D48174 N48174 0 diode
R48175 N48174 N48175 10
D48175 N48175 0 diode
R48176 N48175 N48176 10
D48176 N48176 0 diode
R48177 N48176 N48177 10
D48177 N48177 0 diode
R48178 N48177 N48178 10
D48178 N48178 0 diode
R48179 N48178 N48179 10
D48179 N48179 0 diode
R48180 N48179 N48180 10
D48180 N48180 0 diode
R48181 N48180 N48181 10
D48181 N48181 0 diode
R48182 N48181 N48182 10
D48182 N48182 0 diode
R48183 N48182 N48183 10
D48183 N48183 0 diode
R48184 N48183 N48184 10
D48184 N48184 0 diode
R48185 N48184 N48185 10
D48185 N48185 0 diode
R48186 N48185 N48186 10
D48186 N48186 0 diode
R48187 N48186 N48187 10
D48187 N48187 0 diode
R48188 N48187 N48188 10
D48188 N48188 0 diode
R48189 N48188 N48189 10
D48189 N48189 0 diode
R48190 N48189 N48190 10
D48190 N48190 0 diode
R48191 N48190 N48191 10
D48191 N48191 0 diode
R48192 N48191 N48192 10
D48192 N48192 0 diode
R48193 N48192 N48193 10
D48193 N48193 0 diode
R48194 N48193 N48194 10
D48194 N48194 0 diode
R48195 N48194 N48195 10
D48195 N48195 0 diode
R48196 N48195 N48196 10
D48196 N48196 0 diode
R48197 N48196 N48197 10
D48197 N48197 0 diode
R48198 N48197 N48198 10
D48198 N48198 0 diode
R48199 N48198 N48199 10
D48199 N48199 0 diode
R48200 N48199 N48200 10
D48200 N48200 0 diode
R48201 N48200 N48201 10
D48201 N48201 0 diode
R48202 N48201 N48202 10
D48202 N48202 0 diode
R48203 N48202 N48203 10
D48203 N48203 0 diode
R48204 N48203 N48204 10
D48204 N48204 0 diode
R48205 N48204 N48205 10
D48205 N48205 0 diode
R48206 N48205 N48206 10
D48206 N48206 0 diode
R48207 N48206 N48207 10
D48207 N48207 0 diode
R48208 N48207 N48208 10
D48208 N48208 0 diode
R48209 N48208 N48209 10
D48209 N48209 0 diode
R48210 N48209 N48210 10
D48210 N48210 0 diode
R48211 N48210 N48211 10
D48211 N48211 0 diode
R48212 N48211 N48212 10
D48212 N48212 0 diode
R48213 N48212 N48213 10
D48213 N48213 0 diode
R48214 N48213 N48214 10
D48214 N48214 0 diode
R48215 N48214 N48215 10
D48215 N48215 0 diode
R48216 N48215 N48216 10
D48216 N48216 0 diode
R48217 N48216 N48217 10
D48217 N48217 0 diode
R48218 N48217 N48218 10
D48218 N48218 0 diode
R48219 N48218 N48219 10
D48219 N48219 0 diode
R48220 N48219 N48220 10
D48220 N48220 0 diode
R48221 N48220 N48221 10
D48221 N48221 0 diode
R48222 N48221 N48222 10
D48222 N48222 0 diode
R48223 N48222 N48223 10
D48223 N48223 0 diode
R48224 N48223 N48224 10
D48224 N48224 0 diode
R48225 N48224 N48225 10
D48225 N48225 0 diode
R48226 N48225 N48226 10
D48226 N48226 0 diode
R48227 N48226 N48227 10
D48227 N48227 0 diode
R48228 N48227 N48228 10
D48228 N48228 0 diode
R48229 N48228 N48229 10
D48229 N48229 0 diode
R48230 N48229 N48230 10
D48230 N48230 0 diode
R48231 N48230 N48231 10
D48231 N48231 0 diode
R48232 N48231 N48232 10
D48232 N48232 0 diode
R48233 N48232 N48233 10
D48233 N48233 0 diode
R48234 N48233 N48234 10
D48234 N48234 0 diode
R48235 N48234 N48235 10
D48235 N48235 0 diode
R48236 N48235 N48236 10
D48236 N48236 0 diode
R48237 N48236 N48237 10
D48237 N48237 0 diode
R48238 N48237 N48238 10
D48238 N48238 0 diode
R48239 N48238 N48239 10
D48239 N48239 0 diode
R48240 N48239 N48240 10
D48240 N48240 0 diode
R48241 N48240 N48241 10
D48241 N48241 0 diode
R48242 N48241 N48242 10
D48242 N48242 0 diode
R48243 N48242 N48243 10
D48243 N48243 0 diode
R48244 N48243 N48244 10
D48244 N48244 0 diode
R48245 N48244 N48245 10
D48245 N48245 0 diode
R48246 N48245 N48246 10
D48246 N48246 0 diode
R48247 N48246 N48247 10
D48247 N48247 0 diode
R48248 N48247 N48248 10
D48248 N48248 0 diode
R48249 N48248 N48249 10
D48249 N48249 0 diode
R48250 N48249 N48250 10
D48250 N48250 0 diode
R48251 N48250 N48251 10
D48251 N48251 0 diode
R48252 N48251 N48252 10
D48252 N48252 0 diode
R48253 N48252 N48253 10
D48253 N48253 0 diode
R48254 N48253 N48254 10
D48254 N48254 0 diode
R48255 N48254 N48255 10
D48255 N48255 0 diode
R48256 N48255 N48256 10
D48256 N48256 0 diode
R48257 N48256 N48257 10
D48257 N48257 0 diode
R48258 N48257 N48258 10
D48258 N48258 0 diode
R48259 N48258 N48259 10
D48259 N48259 0 diode
R48260 N48259 N48260 10
D48260 N48260 0 diode
R48261 N48260 N48261 10
D48261 N48261 0 diode
R48262 N48261 N48262 10
D48262 N48262 0 diode
R48263 N48262 N48263 10
D48263 N48263 0 diode
R48264 N48263 N48264 10
D48264 N48264 0 diode
R48265 N48264 N48265 10
D48265 N48265 0 diode
R48266 N48265 N48266 10
D48266 N48266 0 diode
R48267 N48266 N48267 10
D48267 N48267 0 diode
R48268 N48267 N48268 10
D48268 N48268 0 diode
R48269 N48268 N48269 10
D48269 N48269 0 diode
R48270 N48269 N48270 10
D48270 N48270 0 diode
R48271 N48270 N48271 10
D48271 N48271 0 diode
R48272 N48271 N48272 10
D48272 N48272 0 diode
R48273 N48272 N48273 10
D48273 N48273 0 diode
R48274 N48273 N48274 10
D48274 N48274 0 diode
R48275 N48274 N48275 10
D48275 N48275 0 diode
R48276 N48275 N48276 10
D48276 N48276 0 diode
R48277 N48276 N48277 10
D48277 N48277 0 diode
R48278 N48277 N48278 10
D48278 N48278 0 diode
R48279 N48278 N48279 10
D48279 N48279 0 diode
R48280 N48279 N48280 10
D48280 N48280 0 diode
R48281 N48280 N48281 10
D48281 N48281 0 diode
R48282 N48281 N48282 10
D48282 N48282 0 diode
R48283 N48282 N48283 10
D48283 N48283 0 diode
R48284 N48283 N48284 10
D48284 N48284 0 diode
R48285 N48284 N48285 10
D48285 N48285 0 diode
R48286 N48285 N48286 10
D48286 N48286 0 diode
R48287 N48286 N48287 10
D48287 N48287 0 diode
R48288 N48287 N48288 10
D48288 N48288 0 diode
R48289 N48288 N48289 10
D48289 N48289 0 diode
R48290 N48289 N48290 10
D48290 N48290 0 diode
R48291 N48290 N48291 10
D48291 N48291 0 diode
R48292 N48291 N48292 10
D48292 N48292 0 diode
R48293 N48292 N48293 10
D48293 N48293 0 diode
R48294 N48293 N48294 10
D48294 N48294 0 diode
R48295 N48294 N48295 10
D48295 N48295 0 diode
R48296 N48295 N48296 10
D48296 N48296 0 diode
R48297 N48296 N48297 10
D48297 N48297 0 diode
R48298 N48297 N48298 10
D48298 N48298 0 diode
R48299 N48298 N48299 10
D48299 N48299 0 diode
R48300 N48299 N48300 10
D48300 N48300 0 diode
R48301 N48300 N48301 10
D48301 N48301 0 diode
R48302 N48301 N48302 10
D48302 N48302 0 diode
R48303 N48302 N48303 10
D48303 N48303 0 diode
R48304 N48303 N48304 10
D48304 N48304 0 diode
R48305 N48304 N48305 10
D48305 N48305 0 diode
R48306 N48305 N48306 10
D48306 N48306 0 diode
R48307 N48306 N48307 10
D48307 N48307 0 diode
R48308 N48307 N48308 10
D48308 N48308 0 diode
R48309 N48308 N48309 10
D48309 N48309 0 diode
R48310 N48309 N48310 10
D48310 N48310 0 diode
R48311 N48310 N48311 10
D48311 N48311 0 diode
R48312 N48311 N48312 10
D48312 N48312 0 diode
R48313 N48312 N48313 10
D48313 N48313 0 diode
R48314 N48313 N48314 10
D48314 N48314 0 diode
R48315 N48314 N48315 10
D48315 N48315 0 diode
R48316 N48315 N48316 10
D48316 N48316 0 diode
R48317 N48316 N48317 10
D48317 N48317 0 diode
R48318 N48317 N48318 10
D48318 N48318 0 diode
R48319 N48318 N48319 10
D48319 N48319 0 diode
R48320 N48319 N48320 10
D48320 N48320 0 diode
R48321 N48320 N48321 10
D48321 N48321 0 diode
R48322 N48321 N48322 10
D48322 N48322 0 diode
R48323 N48322 N48323 10
D48323 N48323 0 diode
R48324 N48323 N48324 10
D48324 N48324 0 diode
R48325 N48324 N48325 10
D48325 N48325 0 diode
R48326 N48325 N48326 10
D48326 N48326 0 diode
R48327 N48326 N48327 10
D48327 N48327 0 diode
R48328 N48327 N48328 10
D48328 N48328 0 diode
R48329 N48328 N48329 10
D48329 N48329 0 diode
R48330 N48329 N48330 10
D48330 N48330 0 diode
R48331 N48330 N48331 10
D48331 N48331 0 diode
R48332 N48331 N48332 10
D48332 N48332 0 diode
R48333 N48332 N48333 10
D48333 N48333 0 diode
R48334 N48333 N48334 10
D48334 N48334 0 diode
R48335 N48334 N48335 10
D48335 N48335 0 diode
R48336 N48335 N48336 10
D48336 N48336 0 diode
R48337 N48336 N48337 10
D48337 N48337 0 diode
R48338 N48337 N48338 10
D48338 N48338 0 diode
R48339 N48338 N48339 10
D48339 N48339 0 diode
R48340 N48339 N48340 10
D48340 N48340 0 diode
R48341 N48340 N48341 10
D48341 N48341 0 diode
R48342 N48341 N48342 10
D48342 N48342 0 diode
R48343 N48342 N48343 10
D48343 N48343 0 diode
R48344 N48343 N48344 10
D48344 N48344 0 diode
R48345 N48344 N48345 10
D48345 N48345 0 diode
R48346 N48345 N48346 10
D48346 N48346 0 diode
R48347 N48346 N48347 10
D48347 N48347 0 diode
R48348 N48347 N48348 10
D48348 N48348 0 diode
R48349 N48348 N48349 10
D48349 N48349 0 diode
R48350 N48349 N48350 10
D48350 N48350 0 diode
R48351 N48350 N48351 10
D48351 N48351 0 diode
R48352 N48351 N48352 10
D48352 N48352 0 diode
R48353 N48352 N48353 10
D48353 N48353 0 diode
R48354 N48353 N48354 10
D48354 N48354 0 diode
R48355 N48354 N48355 10
D48355 N48355 0 diode
R48356 N48355 N48356 10
D48356 N48356 0 diode
R48357 N48356 N48357 10
D48357 N48357 0 diode
R48358 N48357 N48358 10
D48358 N48358 0 diode
R48359 N48358 N48359 10
D48359 N48359 0 diode
R48360 N48359 N48360 10
D48360 N48360 0 diode
R48361 N48360 N48361 10
D48361 N48361 0 diode
R48362 N48361 N48362 10
D48362 N48362 0 diode
R48363 N48362 N48363 10
D48363 N48363 0 diode
R48364 N48363 N48364 10
D48364 N48364 0 diode
R48365 N48364 N48365 10
D48365 N48365 0 diode
R48366 N48365 N48366 10
D48366 N48366 0 diode
R48367 N48366 N48367 10
D48367 N48367 0 diode
R48368 N48367 N48368 10
D48368 N48368 0 diode
R48369 N48368 N48369 10
D48369 N48369 0 diode
R48370 N48369 N48370 10
D48370 N48370 0 diode
R48371 N48370 N48371 10
D48371 N48371 0 diode
R48372 N48371 N48372 10
D48372 N48372 0 diode
R48373 N48372 N48373 10
D48373 N48373 0 diode
R48374 N48373 N48374 10
D48374 N48374 0 diode
R48375 N48374 N48375 10
D48375 N48375 0 diode
R48376 N48375 N48376 10
D48376 N48376 0 diode
R48377 N48376 N48377 10
D48377 N48377 0 diode
R48378 N48377 N48378 10
D48378 N48378 0 diode
R48379 N48378 N48379 10
D48379 N48379 0 diode
R48380 N48379 N48380 10
D48380 N48380 0 diode
R48381 N48380 N48381 10
D48381 N48381 0 diode
R48382 N48381 N48382 10
D48382 N48382 0 diode
R48383 N48382 N48383 10
D48383 N48383 0 diode
R48384 N48383 N48384 10
D48384 N48384 0 diode
R48385 N48384 N48385 10
D48385 N48385 0 diode
R48386 N48385 N48386 10
D48386 N48386 0 diode
R48387 N48386 N48387 10
D48387 N48387 0 diode
R48388 N48387 N48388 10
D48388 N48388 0 diode
R48389 N48388 N48389 10
D48389 N48389 0 diode
R48390 N48389 N48390 10
D48390 N48390 0 diode
R48391 N48390 N48391 10
D48391 N48391 0 diode
R48392 N48391 N48392 10
D48392 N48392 0 diode
R48393 N48392 N48393 10
D48393 N48393 0 diode
R48394 N48393 N48394 10
D48394 N48394 0 diode
R48395 N48394 N48395 10
D48395 N48395 0 diode
R48396 N48395 N48396 10
D48396 N48396 0 diode
R48397 N48396 N48397 10
D48397 N48397 0 diode
R48398 N48397 N48398 10
D48398 N48398 0 diode
R48399 N48398 N48399 10
D48399 N48399 0 diode
R48400 N48399 N48400 10
D48400 N48400 0 diode
R48401 N48400 N48401 10
D48401 N48401 0 diode
R48402 N48401 N48402 10
D48402 N48402 0 diode
R48403 N48402 N48403 10
D48403 N48403 0 diode
R48404 N48403 N48404 10
D48404 N48404 0 diode
R48405 N48404 N48405 10
D48405 N48405 0 diode
R48406 N48405 N48406 10
D48406 N48406 0 diode
R48407 N48406 N48407 10
D48407 N48407 0 diode
R48408 N48407 N48408 10
D48408 N48408 0 diode
R48409 N48408 N48409 10
D48409 N48409 0 diode
R48410 N48409 N48410 10
D48410 N48410 0 diode
R48411 N48410 N48411 10
D48411 N48411 0 diode
R48412 N48411 N48412 10
D48412 N48412 0 diode
R48413 N48412 N48413 10
D48413 N48413 0 diode
R48414 N48413 N48414 10
D48414 N48414 0 diode
R48415 N48414 N48415 10
D48415 N48415 0 diode
R48416 N48415 N48416 10
D48416 N48416 0 diode
R48417 N48416 N48417 10
D48417 N48417 0 diode
R48418 N48417 N48418 10
D48418 N48418 0 diode
R48419 N48418 N48419 10
D48419 N48419 0 diode
R48420 N48419 N48420 10
D48420 N48420 0 diode
R48421 N48420 N48421 10
D48421 N48421 0 diode
R48422 N48421 N48422 10
D48422 N48422 0 diode
R48423 N48422 N48423 10
D48423 N48423 0 diode
R48424 N48423 N48424 10
D48424 N48424 0 diode
R48425 N48424 N48425 10
D48425 N48425 0 diode
R48426 N48425 N48426 10
D48426 N48426 0 diode
R48427 N48426 N48427 10
D48427 N48427 0 diode
R48428 N48427 N48428 10
D48428 N48428 0 diode
R48429 N48428 N48429 10
D48429 N48429 0 diode
R48430 N48429 N48430 10
D48430 N48430 0 diode
R48431 N48430 N48431 10
D48431 N48431 0 diode
R48432 N48431 N48432 10
D48432 N48432 0 diode
R48433 N48432 N48433 10
D48433 N48433 0 diode
R48434 N48433 N48434 10
D48434 N48434 0 diode
R48435 N48434 N48435 10
D48435 N48435 0 diode
R48436 N48435 N48436 10
D48436 N48436 0 diode
R48437 N48436 N48437 10
D48437 N48437 0 diode
R48438 N48437 N48438 10
D48438 N48438 0 diode
R48439 N48438 N48439 10
D48439 N48439 0 diode
R48440 N48439 N48440 10
D48440 N48440 0 diode
R48441 N48440 N48441 10
D48441 N48441 0 diode
R48442 N48441 N48442 10
D48442 N48442 0 diode
R48443 N48442 N48443 10
D48443 N48443 0 diode
R48444 N48443 N48444 10
D48444 N48444 0 diode
R48445 N48444 N48445 10
D48445 N48445 0 diode
R48446 N48445 N48446 10
D48446 N48446 0 diode
R48447 N48446 N48447 10
D48447 N48447 0 diode
R48448 N48447 N48448 10
D48448 N48448 0 diode
R48449 N48448 N48449 10
D48449 N48449 0 diode
R48450 N48449 N48450 10
D48450 N48450 0 diode
R48451 N48450 N48451 10
D48451 N48451 0 diode
R48452 N48451 N48452 10
D48452 N48452 0 diode
R48453 N48452 N48453 10
D48453 N48453 0 diode
R48454 N48453 N48454 10
D48454 N48454 0 diode
R48455 N48454 N48455 10
D48455 N48455 0 diode
R48456 N48455 N48456 10
D48456 N48456 0 diode
R48457 N48456 N48457 10
D48457 N48457 0 diode
R48458 N48457 N48458 10
D48458 N48458 0 diode
R48459 N48458 N48459 10
D48459 N48459 0 diode
R48460 N48459 N48460 10
D48460 N48460 0 diode
R48461 N48460 N48461 10
D48461 N48461 0 diode
R48462 N48461 N48462 10
D48462 N48462 0 diode
R48463 N48462 N48463 10
D48463 N48463 0 diode
R48464 N48463 N48464 10
D48464 N48464 0 diode
R48465 N48464 N48465 10
D48465 N48465 0 diode
R48466 N48465 N48466 10
D48466 N48466 0 diode
R48467 N48466 N48467 10
D48467 N48467 0 diode
R48468 N48467 N48468 10
D48468 N48468 0 diode
R48469 N48468 N48469 10
D48469 N48469 0 diode
R48470 N48469 N48470 10
D48470 N48470 0 diode
R48471 N48470 N48471 10
D48471 N48471 0 diode
R48472 N48471 N48472 10
D48472 N48472 0 diode
R48473 N48472 N48473 10
D48473 N48473 0 diode
R48474 N48473 N48474 10
D48474 N48474 0 diode
R48475 N48474 N48475 10
D48475 N48475 0 diode
R48476 N48475 N48476 10
D48476 N48476 0 diode
R48477 N48476 N48477 10
D48477 N48477 0 diode
R48478 N48477 N48478 10
D48478 N48478 0 diode
R48479 N48478 N48479 10
D48479 N48479 0 diode
R48480 N48479 N48480 10
D48480 N48480 0 diode
R48481 N48480 N48481 10
D48481 N48481 0 diode
R48482 N48481 N48482 10
D48482 N48482 0 diode
R48483 N48482 N48483 10
D48483 N48483 0 diode
R48484 N48483 N48484 10
D48484 N48484 0 diode
R48485 N48484 N48485 10
D48485 N48485 0 diode
R48486 N48485 N48486 10
D48486 N48486 0 diode
R48487 N48486 N48487 10
D48487 N48487 0 diode
R48488 N48487 N48488 10
D48488 N48488 0 diode
R48489 N48488 N48489 10
D48489 N48489 0 diode
R48490 N48489 N48490 10
D48490 N48490 0 diode
R48491 N48490 N48491 10
D48491 N48491 0 diode
R48492 N48491 N48492 10
D48492 N48492 0 diode
R48493 N48492 N48493 10
D48493 N48493 0 diode
R48494 N48493 N48494 10
D48494 N48494 0 diode
R48495 N48494 N48495 10
D48495 N48495 0 diode
R48496 N48495 N48496 10
D48496 N48496 0 diode
R48497 N48496 N48497 10
D48497 N48497 0 diode
R48498 N48497 N48498 10
D48498 N48498 0 diode
R48499 N48498 N48499 10
D48499 N48499 0 diode
R48500 N48499 N48500 10
D48500 N48500 0 diode
R48501 N48500 N48501 10
D48501 N48501 0 diode
R48502 N48501 N48502 10
D48502 N48502 0 diode
R48503 N48502 N48503 10
D48503 N48503 0 diode
R48504 N48503 N48504 10
D48504 N48504 0 diode
R48505 N48504 N48505 10
D48505 N48505 0 diode
R48506 N48505 N48506 10
D48506 N48506 0 diode
R48507 N48506 N48507 10
D48507 N48507 0 diode
R48508 N48507 N48508 10
D48508 N48508 0 diode
R48509 N48508 N48509 10
D48509 N48509 0 diode
R48510 N48509 N48510 10
D48510 N48510 0 diode
R48511 N48510 N48511 10
D48511 N48511 0 diode
R48512 N48511 N48512 10
D48512 N48512 0 diode
R48513 N48512 N48513 10
D48513 N48513 0 diode
R48514 N48513 N48514 10
D48514 N48514 0 diode
R48515 N48514 N48515 10
D48515 N48515 0 diode
R48516 N48515 N48516 10
D48516 N48516 0 diode
R48517 N48516 N48517 10
D48517 N48517 0 diode
R48518 N48517 N48518 10
D48518 N48518 0 diode
R48519 N48518 N48519 10
D48519 N48519 0 diode
R48520 N48519 N48520 10
D48520 N48520 0 diode
R48521 N48520 N48521 10
D48521 N48521 0 diode
R48522 N48521 N48522 10
D48522 N48522 0 diode
R48523 N48522 N48523 10
D48523 N48523 0 diode
R48524 N48523 N48524 10
D48524 N48524 0 diode
R48525 N48524 N48525 10
D48525 N48525 0 diode
R48526 N48525 N48526 10
D48526 N48526 0 diode
R48527 N48526 N48527 10
D48527 N48527 0 diode
R48528 N48527 N48528 10
D48528 N48528 0 diode
R48529 N48528 N48529 10
D48529 N48529 0 diode
R48530 N48529 N48530 10
D48530 N48530 0 diode
R48531 N48530 N48531 10
D48531 N48531 0 diode
R48532 N48531 N48532 10
D48532 N48532 0 diode
R48533 N48532 N48533 10
D48533 N48533 0 diode
R48534 N48533 N48534 10
D48534 N48534 0 diode
R48535 N48534 N48535 10
D48535 N48535 0 diode
R48536 N48535 N48536 10
D48536 N48536 0 diode
R48537 N48536 N48537 10
D48537 N48537 0 diode
R48538 N48537 N48538 10
D48538 N48538 0 diode
R48539 N48538 N48539 10
D48539 N48539 0 diode
R48540 N48539 N48540 10
D48540 N48540 0 diode
R48541 N48540 N48541 10
D48541 N48541 0 diode
R48542 N48541 N48542 10
D48542 N48542 0 diode
R48543 N48542 N48543 10
D48543 N48543 0 diode
R48544 N48543 N48544 10
D48544 N48544 0 diode
R48545 N48544 N48545 10
D48545 N48545 0 diode
R48546 N48545 N48546 10
D48546 N48546 0 diode
R48547 N48546 N48547 10
D48547 N48547 0 diode
R48548 N48547 N48548 10
D48548 N48548 0 diode
R48549 N48548 N48549 10
D48549 N48549 0 diode
R48550 N48549 N48550 10
D48550 N48550 0 diode
R48551 N48550 N48551 10
D48551 N48551 0 diode
R48552 N48551 N48552 10
D48552 N48552 0 diode
R48553 N48552 N48553 10
D48553 N48553 0 diode
R48554 N48553 N48554 10
D48554 N48554 0 diode
R48555 N48554 N48555 10
D48555 N48555 0 diode
R48556 N48555 N48556 10
D48556 N48556 0 diode
R48557 N48556 N48557 10
D48557 N48557 0 diode
R48558 N48557 N48558 10
D48558 N48558 0 diode
R48559 N48558 N48559 10
D48559 N48559 0 diode
R48560 N48559 N48560 10
D48560 N48560 0 diode
R48561 N48560 N48561 10
D48561 N48561 0 diode
R48562 N48561 N48562 10
D48562 N48562 0 diode
R48563 N48562 N48563 10
D48563 N48563 0 diode
R48564 N48563 N48564 10
D48564 N48564 0 diode
R48565 N48564 N48565 10
D48565 N48565 0 diode
R48566 N48565 N48566 10
D48566 N48566 0 diode
R48567 N48566 N48567 10
D48567 N48567 0 diode
R48568 N48567 N48568 10
D48568 N48568 0 diode
R48569 N48568 N48569 10
D48569 N48569 0 diode
R48570 N48569 N48570 10
D48570 N48570 0 diode
R48571 N48570 N48571 10
D48571 N48571 0 diode
R48572 N48571 N48572 10
D48572 N48572 0 diode
R48573 N48572 N48573 10
D48573 N48573 0 diode
R48574 N48573 N48574 10
D48574 N48574 0 diode
R48575 N48574 N48575 10
D48575 N48575 0 diode
R48576 N48575 N48576 10
D48576 N48576 0 diode
R48577 N48576 N48577 10
D48577 N48577 0 diode
R48578 N48577 N48578 10
D48578 N48578 0 diode
R48579 N48578 N48579 10
D48579 N48579 0 diode
R48580 N48579 N48580 10
D48580 N48580 0 diode
R48581 N48580 N48581 10
D48581 N48581 0 diode
R48582 N48581 N48582 10
D48582 N48582 0 diode
R48583 N48582 N48583 10
D48583 N48583 0 diode
R48584 N48583 N48584 10
D48584 N48584 0 diode
R48585 N48584 N48585 10
D48585 N48585 0 diode
R48586 N48585 N48586 10
D48586 N48586 0 diode
R48587 N48586 N48587 10
D48587 N48587 0 diode
R48588 N48587 N48588 10
D48588 N48588 0 diode
R48589 N48588 N48589 10
D48589 N48589 0 diode
R48590 N48589 N48590 10
D48590 N48590 0 diode
R48591 N48590 N48591 10
D48591 N48591 0 diode
R48592 N48591 N48592 10
D48592 N48592 0 diode
R48593 N48592 N48593 10
D48593 N48593 0 diode
R48594 N48593 N48594 10
D48594 N48594 0 diode
R48595 N48594 N48595 10
D48595 N48595 0 diode
R48596 N48595 N48596 10
D48596 N48596 0 diode
R48597 N48596 N48597 10
D48597 N48597 0 diode
R48598 N48597 N48598 10
D48598 N48598 0 diode
R48599 N48598 N48599 10
D48599 N48599 0 diode
R48600 N48599 N48600 10
D48600 N48600 0 diode
R48601 N48600 N48601 10
D48601 N48601 0 diode
R48602 N48601 N48602 10
D48602 N48602 0 diode
R48603 N48602 N48603 10
D48603 N48603 0 diode
R48604 N48603 N48604 10
D48604 N48604 0 diode
R48605 N48604 N48605 10
D48605 N48605 0 diode
R48606 N48605 N48606 10
D48606 N48606 0 diode
R48607 N48606 N48607 10
D48607 N48607 0 diode
R48608 N48607 N48608 10
D48608 N48608 0 diode
R48609 N48608 N48609 10
D48609 N48609 0 diode
R48610 N48609 N48610 10
D48610 N48610 0 diode
R48611 N48610 N48611 10
D48611 N48611 0 diode
R48612 N48611 N48612 10
D48612 N48612 0 diode
R48613 N48612 N48613 10
D48613 N48613 0 diode
R48614 N48613 N48614 10
D48614 N48614 0 diode
R48615 N48614 N48615 10
D48615 N48615 0 diode
R48616 N48615 N48616 10
D48616 N48616 0 diode
R48617 N48616 N48617 10
D48617 N48617 0 diode
R48618 N48617 N48618 10
D48618 N48618 0 diode
R48619 N48618 N48619 10
D48619 N48619 0 diode
R48620 N48619 N48620 10
D48620 N48620 0 diode
R48621 N48620 N48621 10
D48621 N48621 0 diode
R48622 N48621 N48622 10
D48622 N48622 0 diode
R48623 N48622 N48623 10
D48623 N48623 0 diode
R48624 N48623 N48624 10
D48624 N48624 0 diode
R48625 N48624 N48625 10
D48625 N48625 0 diode
R48626 N48625 N48626 10
D48626 N48626 0 diode
R48627 N48626 N48627 10
D48627 N48627 0 diode
R48628 N48627 N48628 10
D48628 N48628 0 diode
R48629 N48628 N48629 10
D48629 N48629 0 diode
R48630 N48629 N48630 10
D48630 N48630 0 diode
R48631 N48630 N48631 10
D48631 N48631 0 diode
R48632 N48631 N48632 10
D48632 N48632 0 diode
R48633 N48632 N48633 10
D48633 N48633 0 diode
R48634 N48633 N48634 10
D48634 N48634 0 diode
R48635 N48634 N48635 10
D48635 N48635 0 diode
R48636 N48635 N48636 10
D48636 N48636 0 diode
R48637 N48636 N48637 10
D48637 N48637 0 diode
R48638 N48637 N48638 10
D48638 N48638 0 diode
R48639 N48638 N48639 10
D48639 N48639 0 diode
R48640 N48639 N48640 10
D48640 N48640 0 diode
R48641 N48640 N48641 10
D48641 N48641 0 diode
R48642 N48641 N48642 10
D48642 N48642 0 diode
R48643 N48642 N48643 10
D48643 N48643 0 diode
R48644 N48643 N48644 10
D48644 N48644 0 diode
R48645 N48644 N48645 10
D48645 N48645 0 diode
R48646 N48645 N48646 10
D48646 N48646 0 diode
R48647 N48646 N48647 10
D48647 N48647 0 diode
R48648 N48647 N48648 10
D48648 N48648 0 diode
R48649 N48648 N48649 10
D48649 N48649 0 diode
R48650 N48649 N48650 10
D48650 N48650 0 diode
R48651 N48650 N48651 10
D48651 N48651 0 diode
R48652 N48651 N48652 10
D48652 N48652 0 diode
R48653 N48652 N48653 10
D48653 N48653 0 diode
R48654 N48653 N48654 10
D48654 N48654 0 diode
R48655 N48654 N48655 10
D48655 N48655 0 diode
R48656 N48655 N48656 10
D48656 N48656 0 diode
R48657 N48656 N48657 10
D48657 N48657 0 diode
R48658 N48657 N48658 10
D48658 N48658 0 diode
R48659 N48658 N48659 10
D48659 N48659 0 diode
R48660 N48659 N48660 10
D48660 N48660 0 diode
R48661 N48660 N48661 10
D48661 N48661 0 diode
R48662 N48661 N48662 10
D48662 N48662 0 diode
R48663 N48662 N48663 10
D48663 N48663 0 diode
R48664 N48663 N48664 10
D48664 N48664 0 diode
R48665 N48664 N48665 10
D48665 N48665 0 diode
R48666 N48665 N48666 10
D48666 N48666 0 diode
R48667 N48666 N48667 10
D48667 N48667 0 diode
R48668 N48667 N48668 10
D48668 N48668 0 diode
R48669 N48668 N48669 10
D48669 N48669 0 diode
R48670 N48669 N48670 10
D48670 N48670 0 diode
R48671 N48670 N48671 10
D48671 N48671 0 diode
R48672 N48671 N48672 10
D48672 N48672 0 diode
R48673 N48672 N48673 10
D48673 N48673 0 diode
R48674 N48673 N48674 10
D48674 N48674 0 diode
R48675 N48674 N48675 10
D48675 N48675 0 diode
R48676 N48675 N48676 10
D48676 N48676 0 diode
R48677 N48676 N48677 10
D48677 N48677 0 diode
R48678 N48677 N48678 10
D48678 N48678 0 diode
R48679 N48678 N48679 10
D48679 N48679 0 diode
R48680 N48679 N48680 10
D48680 N48680 0 diode
R48681 N48680 N48681 10
D48681 N48681 0 diode
R48682 N48681 N48682 10
D48682 N48682 0 diode
R48683 N48682 N48683 10
D48683 N48683 0 diode
R48684 N48683 N48684 10
D48684 N48684 0 diode
R48685 N48684 N48685 10
D48685 N48685 0 diode
R48686 N48685 N48686 10
D48686 N48686 0 diode
R48687 N48686 N48687 10
D48687 N48687 0 diode
R48688 N48687 N48688 10
D48688 N48688 0 diode
R48689 N48688 N48689 10
D48689 N48689 0 diode
R48690 N48689 N48690 10
D48690 N48690 0 diode
R48691 N48690 N48691 10
D48691 N48691 0 diode
R48692 N48691 N48692 10
D48692 N48692 0 diode
R48693 N48692 N48693 10
D48693 N48693 0 diode
R48694 N48693 N48694 10
D48694 N48694 0 diode
R48695 N48694 N48695 10
D48695 N48695 0 diode
R48696 N48695 N48696 10
D48696 N48696 0 diode
R48697 N48696 N48697 10
D48697 N48697 0 diode
R48698 N48697 N48698 10
D48698 N48698 0 diode
R48699 N48698 N48699 10
D48699 N48699 0 diode
R48700 N48699 N48700 10
D48700 N48700 0 diode
R48701 N48700 N48701 10
D48701 N48701 0 diode
R48702 N48701 N48702 10
D48702 N48702 0 diode
R48703 N48702 N48703 10
D48703 N48703 0 diode
R48704 N48703 N48704 10
D48704 N48704 0 diode
R48705 N48704 N48705 10
D48705 N48705 0 diode
R48706 N48705 N48706 10
D48706 N48706 0 diode
R48707 N48706 N48707 10
D48707 N48707 0 diode
R48708 N48707 N48708 10
D48708 N48708 0 diode
R48709 N48708 N48709 10
D48709 N48709 0 diode
R48710 N48709 N48710 10
D48710 N48710 0 diode
R48711 N48710 N48711 10
D48711 N48711 0 diode
R48712 N48711 N48712 10
D48712 N48712 0 diode
R48713 N48712 N48713 10
D48713 N48713 0 diode
R48714 N48713 N48714 10
D48714 N48714 0 diode
R48715 N48714 N48715 10
D48715 N48715 0 diode
R48716 N48715 N48716 10
D48716 N48716 0 diode
R48717 N48716 N48717 10
D48717 N48717 0 diode
R48718 N48717 N48718 10
D48718 N48718 0 diode
R48719 N48718 N48719 10
D48719 N48719 0 diode
R48720 N48719 N48720 10
D48720 N48720 0 diode
R48721 N48720 N48721 10
D48721 N48721 0 diode
R48722 N48721 N48722 10
D48722 N48722 0 diode
R48723 N48722 N48723 10
D48723 N48723 0 diode
R48724 N48723 N48724 10
D48724 N48724 0 diode
R48725 N48724 N48725 10
D48725 N48725 0 diode
R48726 N48725 N48726 10
D48726 N48726 0 diode
R48727 N48726 N48727 10
D48727 N48727 0 diode
R48728 N48727 N48728 10
D48728 N48728 0 diode
R48729 N48728 N48729 10
D48729 N48729 0 diode
R48730 N48729 N48730 10
D48730 N48730 0 diode
R48731 N48730 N48731 10
D48731 N48731 0 diode
R48732 N48731 N48732 10
D48732 N48732 0 diode
R48733 N48732 N48733 10
D48733 N48733 0 diode
R48734 N48733 N48734 10
D48734 N48734 0 diode
R48735 N48734 N48735 10
D48735 N48735 0 diode
R48736 N48735 N48736 10
D48736 N48736 0 diode
R48737 N48736 N48737 10
D48737 N48737 0 diode
R48738 N48737 N48738 10
D48738 N48738 0 diode
R48739 N48738 N48739 10
D48739 N48739 0 diode
R48740 N48739 N48740 10
D48740 N48740 0 diode
R48741 N48740 N48741 10
D48741 N48741 0 diode
R48742 N48741 N48742 10
D48742 N48742 0 diode
R48743 N48742 N48743 10
D48743 N48743 0 diode
R48744 N48743 N48744 10
D48744 N48744 0 diode
R48745 N48744 N48745 10
D48745 N48745 0 diode
R48746 N48745 N48746 10
D48746 N48746 0 diode
R48747 N48746 N48747 10
D48747 N48747 0 diode
R48748 N48747 N48748 10
D48748 N48748 0 diode
R48749 N48748 N48749 10
D48749 N48749 0 diode
R48750 N48749 N48750 10
D48750 N48750 0 diode
R48751 N48750 N48751 10
D48751 N48751 0 diode
R48752 N48751 N48752 10
D48752 N48752 0 diode
R48753 N48752 N48753 10
D48753 N48753 0 diode
R48754 N48753 N48754 10
D48754 N48754 0 diode
R48755 N48754 N48755 10
D48755 N48755 0 diode
R48756 N48755 N48756 10
D48756 N48756 0 diode
R48757 N48756 N48757 10
D48757 N48757 0 diode
R48758 N48757 N48758 10
D48758 N48758 0 diode
R48759 N48758 N48759 10
D48759 N48759 0 diode
R48760 N48759 N48760 10
D48760 N48760 0 diode
R48761 N48760 N48761 10
D48761 N48761 0 diode
R48762 N48761 N48762 10
D48762 N48762 0 diode
R48763 N48762 N48763 10
D48763 N48763 0 diode
R48764 N48763 N48764 10
D48764 N48764 0 diode
R48765 N48764 N48765 10
D48765 N48765 0 diode
R48766 N48765 N48766 10
D48766 N48766 0 diode
R48767 N48766 N48767 10
D48767 N48767 0 diode
R48768 N48767 N48768 10
D48768 N48768 0 diode
R48769 N48768 N48769 10
D48769 N48769 0 diode
R48770 N48769 N48770 10
D48770 N48770 0 diode
R48771 N48770 N48771 10
D48771 N48771 0 diode
R48772 N48771 N48772 10
D48772 N48772 0 diode
R48773 N48772 N48773 10
D48773 N48773 0 diode
R48774 N48773 N48774 10
D48774 N48774 0 diode
R48775 N48774 N48775 10
D48775 N48775 0 diode
R48776 N48775 N48776 10
D48776 N48776 0 diode
R48777 N48776 N48777 10
D48777 N48777 0 diode
R48778 N48777 N48778 10
D48778 N48778 0 diode
R48779 N48778 N48779 10
D48779 N48779 0 diode
R48780 N48779 N48780 10
D48780 N48780 0 diode
R48781 N48780 N48781 10
D48781 N48781 0 diode
R48782 N48781 N48782 10
D48782 N48782 0 diode
R48783 N48782 N48783 10
D48783 N48783 0 diode
R48784 N48783 N48784 10
D48784 N48784 0 diode
R48785 N48784 N48785 10
D48785 N48785 0 diode
R48786 N48785 N48786 10
D48786 N48786 0 diode
R48787 N48786 N48787 10
D48787 N48787 0 diode
R48788 N48787 N48788 10
D48788 N48788 0 diode
R48789 N48788 N48789 10
D48789 N48789 0 diode
R48790 N48789 N48790 10
D48790 N48790 0 diode
R48791 N48790 N48791 10
D48791 N48791 0 diode
R48792 N48791 N48792 10
D48792 N48792 0 diode
R48793 N48792 N48793 10
D48793 N48793 0 diode
R48794 N48793 N48794 10
D48794 N48794 0 diode
R48795 N48794 N48795 10
D48795 N48795 0 diode
R48796 N48795 N48796 10
D48796 N48796 0 diode
R48797 N48796 N48797 10
D48797 N48797 0 diode
R48798 N48797 N48798 10
D48798 N48798 0 diode
R48799 N48798 N48799 10
D48799 N48799 0 diode
R48800 N48799 N48800 10
D48800 N48800 0 diode
R48801 N48800 N48801 10
D48801 N48801 0 diode
R48802 N48801 N48802 10
D48802 N48802 0 diode
R48803 N48802 N48803 10
D48803 N48803 0 diode
R48804 N48803 N48804 10
D48804 N48804 0 diode
R48805 N48804 N48805 10
D48805 N48805 0 diode
R48806 N48805 N48806 10
D48806 N48806 0 diode
R48807 N48806 N48807 10
D48807 N48807 0 diode
R48808 N48807 N48808 10
D48808 N48808 0 diode
R48809 N48808 N48809 10
D48809 N48809 0 diode
R48810 N48809 N48810 10
D48810 N48810 0 diode
R48811 N48810 N48811 10
D48811 N48811 0 diode
R48812 N48811 N48812 10
D48812 N48812 0 diode
R48813 N48812 N48813 10
D48813 N48813 0 diode
R48814 N48813 N48814 10
D48814 N48814 0 diode
R48815 N48814 N48815 10
D48815 N48815 0 diode
R48816 N48815 N48816 10
D48816 N48816 0 diode
R48817 N48816 N48817 10
D48817 N48817 0 diode
R48818 N48817 N48818 10
D48818 N48818 0 diode
R48819 N48818 N48819 10
D48819 N48819 0 diode
R48820 N48819 N48820 10
D48820 N48820 0 diode
R48821 N48820 N48821 10
D48821 N48821 0 diode
R48822 N48821 N48822 10
D48822 N48822 0 diode
R48823 N48822 N48823 10
D48823 N48823 0 diode
R48824 N48823 N48824 10
D48824 N48824 0 diode
R48825 N48824 N48825 10
D48825 N48825 0 diode
R48826 N48825 N48826 10
D48826 N48826 0 diode
R48827 N48826 N48827 10
D48827 N48827 0 diode
R48828 N48827 N48828 10
D48828 N48828 0 diode
R48829 N48828 N48829 10
D48829 N48829 0 diode
R48830 N48829 N48830 10
D48830 N48830 0 diode
R48831 N48830 N48831 10
D48831 N48831 0 diode
R48832 N48831 N48832 10
D48832 N48832 0 diode
R48833 N48832 N48833 10
D48833 N48833 0 diode
R48834 N48833 N48834 10
D48834 N48834 0 diode
R48835 N48834 N48835 10
D48835 N48835 0 diode
R48836 N48835 N48836 10
D48836 N48836 0 diode
R48837 N48836 N48837 10
D48837 N48837 0 diode
R48838 N48837 N48838 10
D48838 N48838 0 diode
R48839 N48838 N48839 10
D48839 N48839 0 diode
R48840 N48839 N48840 10
D48840 N48840 0 diode
R48841 N48840 N48841 10
D48841 N48841 0 diode
R48842 N48841 N48842 10
D48842 N48842 0 diode
R48843 N48842 N48843 10
D48843 N48843 0 diode
R48844 N48843 N48844 10
D48844 N48844 0 diode
R48845 N48844 N48845 10
D48845 N48845 0 diode
R48846 N48845 N48846 10
D48846 N48846 0 diode
R48847 N48846 N48847 10
D48847 N48847 0 diode
R48848 N48847 N48848 10
D48848 N48848 0 diode
R48849 N48848 N48849 10
D48849 N48849 0 diode
R48850 N48849 N48850 10
D48850 N48850 0 diode
R48851 N48850 N48851 10
D48851 N48851 0 diode
R48852 N48851 N48852 10
D48852 N48852 0 diode
R48853 N48852 N48853 10
D48853 N48853 0 diode
R48854 N48853 N48854 10
D48854 N48854 0 diode
R48855 N48854 N48855 10
D48855 N48855 0 diode
R48856 N48855 N48856 10
D48856 N48856 0 diode
R48857 N48856 N48857 10
D48857 N48857 0 diode
R48858 N48857 N48858 10
D48858 N48858 0 diode
R48859 N48858 N48859 10
D48859 N48859 0 diode
R48860 N48859 N48860 10
D48860 N48860 0 diode
R48861 N48860 N48861 10
D48861 N48861 0 diode
R48862 N48861 N48862 10
D48862 N48862 0 diode
R48863 N48862 N48863 10
D48863 N48863 0 diode
R48864 N48863 N48864 10
D48864 N48864 0 diode
R48865 N48864 N48865 10
D48865 N48865 0 diode
R48866 N48865 N48866 10
D48866 N48866 0 diode
R48867 N48866 N48867 10
D48867 N48867 0 diode
R48868 N48867 N48868 10
D48868 N48868 0 diode
R48869 N48868 N48869 10
D48869 N48869 0 diode
R48870 N48869 N48870 10
D48870 N48870 0 diode
R48871 N48870 N48871 10
D48871 N48871 0 diode
R48872 N48871 N48872 10
D48872 N48872 0 diode
R48873 N48872 N48873 10
D48873 N48873 0 diode
R48874 N48873 N48874 10
D48874 N48874 0 diode
R48875 N48874 N48875 10
D48875 N48875 0 diode
R48876 N48875 N48876 10
D48876 N48876 0 diode
R48877 N48876 N48877 10
D48877 N48877 0 diode
R48878 N48877 N48878 10
D48878 N48878 0 diode
R48879 N48878 N48879 10
D48879 N48879 0 diode
R48880 N48879 N48880 10
D48880 N48880 0 diode
R48881 N48880 N48881 10
D48881 N48881 0 diode
R48882 N48881 N48882 10
D48882 N48882 0 diode
R48883 N48882 N48883 10
D48883 N48883 0 diode
R48884 N48883 N48884 10
D48884 N48884 0 diode
R48885 N48884 N48885 10
D48885 N48885 0 diode
R48886 N48885 N48886 10
D48886 N48886 0 diode
R48887 N48886 N48887 10
D48887 N48887 0 diode
R48888 N48887 N48888 10
D48888 N48888 0 diode
R48889 N48888 N48889 10
D48889 N48889 0 diode
R48890 N48889 N48890 10
D48890 N48890 0 diode
R48891 N48890 N48891 10
D48891 N48891 0 diode
R48892 N48891 N48892 10
D48892 N48892 0 diode
R48893 N48892 N48893 10
D48893 N48893 0 diode
R48894 N48893 N48894 10
D48894 N48894 0 diode
R48895 N48894 N48895 10
D48895 N48895 0 diode
R48896 N48895 N48896 10
D48896 N48896 0 diode
R48897 N48896 N48897 10
D48897 N48897 0 diode
R48898 N48897 N48898 10
D48898 N48898 0 diode
R48899 N48898 N48899 10
D48899 N48899 0 diode
R48900 N48899 N48900 10
D48900 N48900 0 diode
R48901 N48900 N48901 10
D48901 N48901 0 diode
R48902 N48901 N48902 10
D48902 N48902 0 diode
R48903 N48902 N48903 10
D48903 N48903 0 diode
R48904 N48903 N48904 10
D48904 N48904 0 diode
R48905 N48904 N48905 10
D48905 N48905 0 diode
R48906 N48905 N48906 10
D48906 N48906 0 diode
R48907 N48906 N48907 10
D48907 N48907 0 diode
R48908 N48907 N48908 10
D48908 N48908 0 diode
R48909 N48908 N48909 10
D48909 N48909 0 diode
R48910 N48909 N48910 10
D48910 N48910 0 diode
R48911 N48910 N48911 10
D48911 N48911 0 diode
R48912 N48911 N48912 10
D48912 N48912 0 diode
R48913 N48912 N48913 10
D48913 N48913 0 diode
R48914 N48913 N48914 10
D48914 N48914 0 diode
R48915 N48914 N48915 10
D48915 N48915 0 diode
R48916 N48915 N48916 10
D48916 N48916 0 diode
R48917 N48916 N48917 10
D48917 N48917 0 diode
R48918 N48917 N48918 10
D48918 N48918 0 diode
R48919 N48918 N48919 10
D48919 N48919 0 diode
R48920 N48919 N48920 10
D48920 N48920 0 diode
R48921 N48920 N48921 10
D48921 N48921 0 diode
R48922 N48921 N48922 10
D48922 N48922 0 diode
R48923 N48922 N48923 10
D48923 N48923 0 diode
R48924 N48923 N48924 10
D48924 N48924 0 diode
R48925 N48924 N48925 10
D48925 N48925 0 diode
R48926 N48925 N48926 10
D48926 N48926 0 diode
R48927 N48926 N48927 10
D48927 N48927 0 diode
R48928 N48927 N48928 10
D48928 N48928 0 diode
R48929 N48928 N48929 10
D48929 N48929 0 diode
R48930 N48929 N48930 10
D48930 N48930 0 diode
R48931 N48930 N48931 10
D48931 N48931 0 diode
R48932 N48931 N48932 10
D48932 N48932 0 diode
R48933 N48932 N48933 10
D48933 N48933 0 diode
R48934 N48933 N48934 10
D48934 N48934 0 diode
R48935 N48934 N48935 10
D48935 N48935 0 diode
R48936 N48935 N48936 10
D48936 N48936 0 diode
R48937 N48936 N48937 10
D48937 N48937 0 diode
R48938 N48937 N48938 10
D48938 N48938 0 diode
R48939 N48938 N48939 10
D48939 N48939 0 diode
R48940 N48939 N48940 10
D48940 N48940 0 diode
R48941 N48940 N48941 10
D48941 N48941 0 diode
R48942 N48941 N48942 10
D48942 N48942 0 diode
R48943 N48942 N48943 10
D48943 N48943 0 diode
R48944 N48943 N48944 10
D48944 N48944 0 diode
R48945 N48944 N48945 10
D48945 N48945 0 diode
R48946 N48945 N48946 10
D48946 N48946 0 diode
R48947 N48946 N48947 10
D48947 N48947 0 diode
R48948 N48947 N48948 10
D48948 N48948 0 diode
R48949 N48948 N48949 10
D48949 N48949 0 diode
R48950 N48949 N48950 10
D48950 N48950 0 diode
R48951 N48950 N48951 10
D48951 N48951 0 diode
R48952 N48951 N48952 10
D48952 N48952 0 diode
R48953 N48952 N48953 10
D48953 N48953 0 diode
R48954 N48953 N48954 10
D48954 N48954 0 diode
R48955 N48954 N48955 10
D48955 N48955 0 diode
R48956 N48955 N48956 10
D48956 N48956 0 diode
R48957 N48956 N48957 10
D48957 N48957 0 diode
R48958 N48957 N48958 10
D48958 N48958 0 diode
R48959 N48958 N48959 10
D48959 N48959 0 diode
R48960 N48959 N48960 10
D48960 N48960 0 diode
R48961 N48960 N48961 10
D48961 N48961 0 diode
R48962 N48961 N48962 10
D48962 N48962 0 diode
R48963 N48962 N48963 10
D48963 N48963 0 diode
R48964 N48963 N48964 10
D48964 N48964 0 diode
R48965 N48964 N48965 10
D48965 N48965 0 diode
R48966 N48965 N48966 10
D48966 N48966 0 diode
R48967 N48966 N48967 10
D48967 N48967 0 diode
R48968 N48967 N48968 10
D48968 N48968 0 diode
R48969 N48968 N48969 10
D48969 N48969 0 diode
R48970 N48969 N48970 10
D48970 N48970 0 diode
R48971 N48970 N48971 10
D48971 N48971 0 diode
R48972 N48971 N48972 10
D48972 N48972 0 diode
R48973 N48972 N48973 10
D48973 N48973 0 diode
R48974 N48973 N48974 10
D48974 N48974 0 diode
R48975 N48974 N48975 10
D48975 N48975 0 diode
R48976 N48975 N48976 10
D48976 N48976 0 diode
R48977 N48976 N48977 10
D48977 N48977 0 diode
R48978 N48977 N48978 10
D48978 N48978 0 diode
R48979 N48978 N48979 10
D48979 N48979 0 diode
R48980 N48979 N48980 10
D48980 N48980 0 diode
R48981 N48980 N48981 10
D48981 N48981 0 diode
R48982 N48981 N48982 10
D48982 N48982 0 diode
R48983 N48982 N48983 10
D48983 N48983 0 diode
R48984 N48983 N48984 10
D48984 N48984 0 diode
R48985 N48984 N48985 10
D48985 N48985 0 diode
R48986 N48985 N48986 10
D48986 N48986 0 diode
R48987 N48986 N48987 10
D48987 N48987 0 diode
R48988 N48987 N48988 10
D48988 N48988 0 diode
R48989 N48988 N48989 10
D48989 N48989 0 diode
R48990 N48989 N48990 10
D48990 N48990 0 diode
R48991 N48990 N48991 10
D48991 N48991 0 diode
R48992 N48991 N48992 10
D48992 N48992 0 diode
R48993 N48992 N48993 10
D48993 N48993 0 diode
R48994 N48993 N48994 10
D48994 N48994 0 diode
R48995 N48994 N48995 10
D48995 N48995 0 diode
R48996 N48995 N48996 10
D48996 N48996 0 diode
R48997 N48996 N48997 10
D48997 N48997 0 diode
R48998 N48997 N48998 10
D48998 N48998 0 diode
R48999 N48998 N48999 10
D48999 N48999 0 diode
R49000 N48999 N49000 10
D49000 N49000 0 diode
R49001 N49000 N49001 10
D49001 N49001 0 diode
R49002 N49001 N49002 10
D49002 N49002 0 diode
R49003 N49002 N49003 10
D49003 N49003 0 diode
R49004 N49003 N49004 10
D49004 N49004 0 diode
R49005 N49004 N49005 10
D49005 N49005 0 diode
R49006 N49005 N49006 10
D49006 N49006 0 diode
R49007 N49006 N49007 10
D49007 N49007 0 diode
R49008 N49007 N49008 10
D49008 N49008 0 diode
R49009 N49008 N49009 10
D49009 N49009 0 diode
R49010 N49009 N49010 10
D49010 N49010 0 diode
R49011 N49010 N49011 10
D49011 N49011 0 diode
R49012 N49011 N49012 10
D49012 N49012 0 diode
R49013 N49012 N49013 10
D49013 N49013 0 diode
R49014 N49013 N49014 10
D49014 N49014 0 diode
R49015 N49014 N49015 10
D49015 N49015 0 diode
R49016 N49015 N49016 10
D49016 N49016 0 diode
R49017 N49016 N49017 10
D49017 N49017 0 diode
R49018 N49017 N49018 10
D49018 N49018 0 diode
R49019 N49018 N49019 10
D49019 N49019 0 diode
R49020 N49019 N49020 10
D49020 N49020 0 diode
R49021 N49020 N49021 10
D49021 N49021 0 diode
R49022 N49021 N49022 10
D49022 N49022 0 diode
R49023 N49022 N49023 10
D49023 N49023 0 diode
R49024 N49023 N49024 10
D49024 N49024 0 diode
R49025 N49024 N49025 10
D49025 N49025 0 diode
R49026 N49025 N49026 10
D49026 N49026 0 diode
R49027 N49026 N49027 10
D49027 N49027 0 diode
R49028 N49027 N49028 10
D49028 N49028 0 diode
R49029 N49028 N49029 10
D49029 N49029 0 diode
R49030 N49029 N49030 10
D49030 N49030 0 diode
R49031 N49030 N49031 10
D49031 N49031 0 diode
R49032 N49031 N49032 10
D49032 N49032 0 diode
R49033 N49032 N49033 10
D49033 N49033 0 diode
R49034 N49033 N49034 10
D49034 N49034 0 diode
R49035 N49034 N49035 10
D49035 N49035 0 diode
R49036 N49035 N49036 10
D49036 N49036 0 diode
R49037 N49036 N49037 10
D49037 N49037 0 diode
R49038 N49037 N49038 10
D49038 N49038 0 diode
R49039 N49038 N49039 10
D49039 N49039 0 diode
R49040 N49039 N49040 10
D49040 N49040 0 diode
R49041 N49040 N49041 10
D49041 N49041 0 diode
R49042 N49041 N49042 10
D49042 N49042 0 diode
R49043 N49042 N49043 10
D49043 N49043 0 diode
R49044 N49043 N49044 10
D49044 N49044 0 diode
R49045 N49044 N49045 10
D49045 N49045 0 diode
R49046 N49045 N49046 10
D49046 N49046 0 diode
R49047 N49046 N49047 10
D49047 N49047 0 diode
R49048 N49047 N49048 10
D49048 N49048 0 diode
R49049 N49048 N49049 10
D49049 N49049 0 diode
R49050 N49049 N49050 10
D49050 N49050 0 diode
R49051 N49050 N49051 10
D49051 N49051 0 diode
R49052 N49051 N49052 10
D49052 N49052 0 diode
R49053 N49052 N49053 10
D49053 N49053 0 diode
R49054 N49053 N49054 10
D49054 N49054 0 diode
R49055 N49054 N49055 10
D49055 N49055 0 diode
R49056 N49055 N49056 10
D49056 N49056 0 diode
R49057 N49056 N49057 10
D49057 N49057 0 diode
R49058 N49057 N49058 10
D49058 N49058 0 diode
R49059 N49058 N49059 10
D49059 N49059 0 diode
R49060 N49059 N49060 10
D49060 N49060 0 diode
R49061 N49060 N49061 10
D49061 N49061 0 diode
R49062 N49061 N49062 10
D49062 N49062 0 diode
R49063 N49062 N49063 10
D49063 N49063 0 diode
R49064 N49063 N49064 10
D49064 N49064 0 diode
R49065 N49064 N49065 10
D49065 N49065 0 diode
R49066 N49065 N49066 10
D49066 N49066 0 diode
R49067 N49066 N49067 10
D49067 N49067 0 diode
R49068 N49067 N49068 10
D49068 N49068 0 diode
R49069 N49068 N49069 10
D49069 N49069 0 diode
R49070 N49069 N49070 10
D49070 N49070 0 diode
R49071 N49070 N49071 10
D49071 N49071 0 diode
R49072 N49071 N49072 10
D49072 N49072 0 diode
R49073 N49072 N49073 10
D49073 N49073 0 diode
R49074 N49073 N49074 10
D49074 N49074 0 diode
R49075 N49074 N49075 10
D49075 N49075 0 diode
R49076 N49075 N49076 10
D49076 N49076 0 diode
R49077 N49076 N49077 10
D49077 N49077 0 diode
R49078 N49077 N49078 10
D49078 N49078 0 diode
R49079 N49078 N49079 10
D49079 N49079 0 diode
R49080 N49079 N49080 10
D49080 N49080 0 diode
R49081 N49080 N49081 10
D49081 N49081 0 diode
R49082 N49081 N49082 10
D49082 N49082 0 diode
R49083 N49082 N49083 10
D49083 N49083 0 diode
R49084 N49083 N49084 10
D49084 N49084 0 diode
R49085 N49084 N49085 10
D49085 N49085 0 diode
R49086 N49085 N49086 10
D49086 N49086 0 diode
R49087 N49086 N49087 10
D49087 N49087 0 diode
R49088 N49087 N49088 10
D49088 N49088 0 diode
R49089 N49088 N49089 10
D49089 N49089 0 diode
R49090 N49089 N49090 10
D49090 N49090 0 diode
R49091 N49090 N49091 10
D49091 N49091 0 diode
R49092 N49091 N49092 10
D49092 N49092 0 diode
R49093 N49092 N49093 10
D49093 N49093 0 diode
R49094 N49093 N49094 10
D49094 N49094 0 diode
R49095 N49094 N49095 10
D49095 N49095 0 diode
R49096 N49095 N49096 10
D49096 N49096 0 diode
R49097 N49096 N49097 10
D49097 N49097 0 diode
R49098 N49097 N49098 10
D49098 N49098 0 diode
R49099 N49098 N49099 10
D49099 N49099 0 diode
R49100 N49099 N49100 10
D49100 N49100 0 diode
R49101 N49100 N49101 10
D49101 N49101 0 diode
R49102 N49101 N49102 10
D49102 N49102 0 diode
R49103 N49102 N49103 10
D49103 N49103 0 diode
R49104 N49103 N49104 10
D49104 N49104 0 diode
R49105 N49104 N49105 10
D49105 N49105 0 diode
R49106 N49105 N49106 10
D49106 N49106 0 diode
R49107 N49106 N49107 10
D49107 N49107 0 diode
R49108 N49107 N49108 10
D49108 N49108 0 diode
R49109 N49108 N49109 10
D49109 N49109 0 diode
R49110 N49109 N49110 10
D49110 N49110 0 diode
R49111 N49110 N49111 10
D49111 N49111 0 diode
R49112 N49111 N49112 10
D49112 N49112 0 diode
R49113 N49112 N49113 10
D49113 N49113 0 diode
R49114 N49113 N49114 10
D49114 N49114 0 diode
R49115 N49114 N49115 10
D49115 N49115 0 diode
R49116 N49115 N49116 10
D49116 N49116 0 diode
R49117 N49116 N49117 10
D49117 N49117 0 diode
R49118 N49117 N49118 10
D49118 N49118 0 diode
R49119 N49118 N49119 10
D49119 N49119 0 diode
R49120 N49119 N49120 10
D49120 N49120 0 diode
R49121 N49120 N49121 10
D49121 N49121 0 diode
R49122 N49121 N49122 10
D49122 N49122 0 diode
R49123 N49122 N49123 10
D49123 N49123 0 diode
R49124 N49123 N49124 10
D49124 N49124 0 diode
R49125 N49124 N49125 10
D49125 N49125 0 diode
R49126 N49125 N49126 10
D49126 N49126 0 diode
R49127 N49126 N49127 10
D49127 N49127 0 diode
R49128 N49127 N49128 10
D49128 N49128 0 diode
R49129 N49128 N49129 10
D49129 N49129 0 diode
R49130 N49129 N49130 10
D49130 N49130 0 diode
R49131 N49130 N49131 10
D49131 N49131 0 diode
R49132 N49131 N49132 10
D49132 N49132 0 diode
R49133 N49132 N49133 10
D49133 N49133 0 diode
R49134 N49133 N49134 10
D49134 N49134 0 diode
R49135 N49134 N49135 10
D49135 N49135 0 diode
R49136 N49135 N49136 10
D49136 N49136 0 diode
R49137 N49136 N49137 10
D49137 N49137 0 diode
R49138 N49137 N49138 10
D49138 N49138 0 diode
R49139 N49138 N49139 10
D49139 N49139 0 diode
R49140 N49139 N49140 10
D49140 N49140 0 diode
R49141 N49140 N49141 10
D49141 N49141 0 diode
R49142 N49141 N49142 10
D49142 N49142 0 diode
R49143 N49142 N49143 10
D49143 N49143 0 diode
R49144 N49143 N49144 10
D49144 N49144 0 diode
R49145 N49144 N49145 10
D49145 N49145 0 diode
R49146 N49145 N49146 10
D49146 N49146 0 diode
R49147 N49146 N49147 10
D49147 N49147 0 diode
R49148 N49147 N49148 10
D49148 N49148 0 diode
R49149 N49148 N49149 10
D49149 N49149 0 diode
R49150 N49149 N49150 10
D49150 N49150 0 diode
R49151 N49150 N49151 10
D49151 N49151 0 diode
R49152 N49151 N49152 10
D49152 N49152 0 diode
R49153 N49152 N49153 10
D49153 N49153 0 diode
R49154 N49153 N49154 10
D49154 N49154 0 diode
R49155 N49154 N49155 10
D49155 N49155 0 diode
R49156 N49155 N49156 10
D49156 N49156 0 diode
R49157 N49156 N49157 10
D49157 N49157 0 diode
R49158 N49157 N49158 10
D49158 N49158 0 diode
R49159 N49158 N49159 10
D49159 N49159 0 diode
R49160 N49159 N49160 10
D49160 N49160 0 diode
R49161 N49160 N49161 10
D49161 N49161 0 diode
R49162 N49161 N49162 10
D49162 N49162 0 diode
R49163 N49162 N49163 10
D49163 N49163 0 diode
R49164 N49163 N49164 10
D49164 N49164 0 diode
R49165 N49164 N49165 10
D49165 N49165 0 diode
R49166 N49165 N49166 10
D49166 N49166 0 diode
R49167 N49166 N49167 10
D49167 N49167 0 diode
R49168 N49167 N49168 10
D49168 N49168 0 diode
R49169 N49168 N49169 10
D49169 N49169 0 diode
R49170 N49169 N49170 10
D49170 N49170 0 diode
R49171 N49170 N49171 10
D49171 N49171 0 diode
R49172 N49171 N49172 10
D49172 N49172 0 diode
R49173 N49172 N49173 10
D49173 N49173 0 diode
R49174 N49173 N49174 10
D49174 N49174 0 diode
R49175 N49174 N49175 10
D49175 N49175 0 diode
R49176 N49175 N49176 10
D49176 N49176 0 diode
R49177 N49176 N49177 10
D49177 N49177 0 diode
R49178 N49177 N49178 10
D49178 N49178 0 diode
R49179 N49178 N49179 10
D49179 N49179 0 diode
R49180 N49179 N49180 10
D49180 N49180 0 diode
R49181 N49180 N49181 10
D49181 N49181 0 diode
R49182 N49181 N49182 10
D49182 N49182 0 diode
R49183 N49182 N49183 10
D49183 N49183 0 diode
R49184 N49183 N49184 10
D49184 N49184 0 diode
R49185 N49184 N49185 10
D49185 N49185 0 diode
R49186 N49185 N49186 10
D49186 N49186 0 diode
R49187 N49186 N49187 10
D49187 N49187 0 diode
R49188 N49187 N49188 10
D49188 N49188 0 diode
R49189 N49188 N49189 10
D49189 N49189 0 diode
R49190 N49189 N49190 10
D49190 N49190 0 diode
R49191 N49190 N49191 10
D49191 N49191 0 diode
R49192 N49191 N49192 10
D49192 N49192 0 diode
R49193 N49192 N49193 10
D49193 N49193 0 diode
R49194 N49193 N49194 10
D49194 N49194 0 diode
R49195 N49194 N49195 10
D49195 N49195 0 diode
R49196 N49195 N49196 10
D49196 N49196 0 diode
R49197 N49196 N49197 10
D49197 N49197 0 diode
R49198 N49197 N49198 10
D49198 N49198 0 diode
R49199 N49198 N49199 10
D49199 N49199 0 diode
R49200 N49199 N49200 10
D49200 N49200 0 diode
R49201 N49200 N49201 10
D49201 N49201 0 diode
R49202 N49201 N49202 10
D49202 N49202 0 diode
R49203 N49202 N49203 10
D49203 N49203 0 diode
R49204 N49203 N49204 10
D49204 N49204 0 diode
R49205 N49204 N49205 10
D49205 N49205 0 diode
R49206 N49205 N49206 10
D49206 N49206 0 diode
R49207 N49206 N49207 10
D49207 N49207 0 diode
R49208 N49207 N49208 10
D49208 N49208 0 diode
R49209 N49208 N49209 10
D49209 N49209 0 diode
R49210 N49209 N49210 10
D49210 N49210 0 diode
R49211 N49210 N49211 10
D49211 N49211 0 diode
R49212 N49211 N49212 10
D49212 N49212 0 diode
R49213 N49212 N49213 10
D49213 N49213 0 diode
R49214 N49213 N49214 10
D49214 N49214 0 diode
R49215 N49214 N49215 10
D49215 N49215 0 diode
R49216 N49215 N49216 10
D49216 N49216 0 diode
R49217 N49216 N49217 10
D49217 N49217 0 diode
R49218 N49217 N49218 10
D49218 N49218 0 diode
R49219 N49218 N49219 10
D49219 N49219 0 diode
R49220 N49219 N49220 10
D49220 N49220 0 diode
R49221 N49220 N49221 10
D49221 N49221 0 diode
R49222 N49221 N49222 10
D49222 N49222 0 diode
R49223 N49222 N49223 10
D49223 N49223 0 diode
R49224 N49223 N49224 10
D49224 N49224 0 diode
R49225 N49224 N49225 10
D49225 N49225 0 diode
R49226 N49225 N49226 10
D49226 N49226 0 diode
R49227 N49226 N49227 10
D49227 N49227 0 diode
R49228 N49227 N49228 10
D49228 N49228 0 diode
R49229 N49228 N49229 10
D49229 N49229 0 diode
R49230 N49229 N49230 10
D49230 N49230 0 diode
R49231 N49230 N49231 10
D49231 N49231 0 diode
R49232 N49231 N49232 10
D49232 N49232 0 diode
R49233 N49232 N49233 10
D49233 N49233 0 diode
R49234 N49233 N49234 10
D49234 N49234 0 diode
R49235 N49234 N49235 10
D49235 N49235 0 diode
R49236 N49235 N49236 10
D49236 N49236 0 diode
R49237 N49236 N49237 10
D49237 N49237 0 diode
R49238 N49237 N49238 10
D49238 N49238 0 diode
R49239 N49238 N49239 10
D49239 N49239 0 diode
R49240 N49239 N49240 10
D49240 N49240 0 diode
R49241 N49240 N49241 10
D49241 N49241 0 diode
R49242 N49241 N49242 10
D49242 N49242 0 diode
R49243 N49242 N49243 10
D49243 N49243 0 diode
R49244 N49243 N49244 10
D49244 N49244 0 diode
R49245 N49244 N49245 10
D49245 N49245 0 diode
R49246 N49245 N49246 10
D49246 N49246 0 diode
R49247 N49246 N49247 10
D49247 N49247 0 diode
R49248 N49247 N49248 10
D49248 N49248 0 diode
R49249 N49248 N49249 10
D49249 N49249 0 diode
R49250 N49249 N49250 10
D49250 N49250 0 diode
R49251 N49250 N49251 10
D49251 N49251 0 diode
R49252 N49251 N49252 10
D49252 N49252 0 diode
R49253 N49252 N49253 10
D49253 N49253 0 diode
R49254 N49253 N49254 10
D49254 N49254 0 diode
R49255 N49254 N49255 10
D49255 N49255 0 diode
R49256 N49255 N49256 10
D49256 N49256 0 diode
R49257 N49256 N49257 10
D49257 N49257 0 diode
R49258 N49257 N49258 10
D49258 N49258 0 diode
R49259 N49258 N49259 10
D49259 N49259 0 diode
R49260 N49259 N49260 10
D49260 N49260 0 diode
R49261 N49260 N49261 10
D49261 N49261 0 diode
R49262 N49261 N49262 10
D49262 N49262 0 diode
R49263 N49262 N49263 10
D49263 N49263 0 diode
R49264 N49263 N49264 10
D49264 N49264 0 diode
R49265 N49264 N49265 10
D49265 N49265 0 diode
R49266 N49265 N49266 10
D49266 N49266 0 diode
R49267 N49266 N49267 10
D49267 N49267 0 diode
R49268 N49267 N49268 10
D49268 N49268 0 diode
R49269 N49268 N49269 10
D49269 N49269 0 diode
R49270 N49269 N49270 10
D49270 N49270 0 diode
R49271 N49270 N49271 10
D49271 N49271 0 diode
R49272 N49271 N49272 10
D49272 N49272 0 diode
R49273 N49272 N49273 10
D49273 N49273 0 diode
R49274 N49273 N49274 10
D49274 N49274 0 diode
R49275 N49274 N49275 10
D49275 N49275 0 diode
R49276 N49275 N49276 10
D49276 N49276 0 diode
R49277 N49276 N49277 10
D49277 N49277 0 diode
R49278 N49277 N49278 10
D49278 N49278 0 diode
R49279 N49278 N49279 10
D49279 N49279 0 diode
R49280 N49279 N49280 10
D49280 N49280 0 diode
R49281 N49280 N49281 10
D49281 N49281 0 diode
R49282 N49281 N49282 10
D49282 N49282 0 diode
R49283 N49282 N49283 10
D49283 N49283 0 diode
R49284 N49283 N49284 10
D49284 N49284 0 diode
R49285 N49284 N49285 10
D49285 N49285 0 diode
R49286 N49285 N49286 10
D49286 N49286 0 diode
R49287 N49286 N49287 10
D49287 N49287 0 diode
R49288 N49287 N49288 10
D49288 N49288 0 diode
R49289 N49288 N49289 10
D49289 N49289 0 diode
R49290 N49289 N49290 10
D49290 N49290 0 diode
R49291 N49290 N49291 10
D49291 N49291 0 diode
R49292 N49291 N49292 10
D49292 N49292 0 diode
R49293 N49292 N49293 10
D49293 N49293 0 diode
R49294 N49293 N49294 10
D49294 N49294 0 diode
R49295 N49294 N49295 10
D49295 N49295 0 diode
R49296 N49295 N49296 10
D49296 N49296 0 diode
R49297 N49296 N49297 10
D49297 N49297 0 diode
R49298 N49297 N49298 10
D49298 N49298 0 diode
R49299 N49298 N49299 10
D49299 N49299 0 diode
R49300 N49299 N49300 10
D49300 N49300 0 diode
R49301 N49300 N49301 10
D49301 N49301 0 diode
R49302 N49301 N49302 10
D49302 N49302 0 diode
R49303 N49302 N49303 10
D49303 N49303 0 diode
R49304 N49303 N49304 10
D49304 N49304 0 diode
R49305 N49304 N49305 10
D49305 N49305 0 diode
R49306 N49305 N49306 10
D49306 N49306 0 diode
R49307 N49306 N49307 10
D49307 N49307 0 diode
R49308 N49307 N49308 10
D49308 N49308 0 diode
R49309 N49308 N49309 10
D49309 N49309 0 diode
R49310 N49309 N49310 10
D49310 N49310 0 diode
R49311 N49310 N49311 10
D49311 N49311 0 diode
R49312 N49311 N49312 10
D49312 N49312 0 diode
R49313 N49312 N49313 10
D49313 N49313 0 diode
R49314 N49313 N49314 10
D49314 N49314 0 diode
R49315 N49314 N49315 10
D49315 N49315 0 diode
R49316 N49315 N49316 10
D49316 N49316 0 diode
R49317 N49316 N49317 10
D49317 N49317 0 diode
R49318 N49317 N49318 10
D49318 N49318 0 diode
R49319 N49318 N49319 10
D49319 N49319 0 diode
R49320 N49319 N49320 10
D49320 N49320 0 diode
R49321 N49320 N49321 10
D49321 N49321 0 diode
R49322 N49321 N49322 10
D49322 N49322 0 diode
R49323 N49322 N49323 10
D49323 N49323 0 diode
R49324 N49323 N49324 10
D49324 N49324 0 diode
R49325 N49324 N49325 10
D49325 N49325 0 diode
R49326 N49325 N49326 10
D49326 N49326 0 diode
R49327 N49326 N49327 10
D49327 N49327 0 diode
R49328 N49327 N49328 10
D49328 N49328 0 diode
R49329 N49328 N49329 10
D49329 N49329 0 diode
R49330 N49329 N49330 10
D49330 N49330 0 diode
R49331 N49330 N49331 10
D49331 N49331 0 diode
R49332 N49331 N49332 10
D49332 N49332 0 diode
R49333 N49332 N49333 10
D49333 N49333 0 diode
R49334 N49333 N49334 10
D49334 N49334 0 diode
R49335 N49334 N49335 10
D49335 N49335 0 diode
R49336 N49335 N49336 10
D49336 N49336 0 diode
R49337 N49336 N49337 10
D49337 N49337 0 diode
R49338 N49337 N49338 10
D49338 N49338 0 diode
R49339 N49338 N49339 10
D49339 N49339 0 diode
R49340 N49339 N49340 10
D49340 N49340 0 diode
R49341 N49340 N49341 10
D49341 N49341 0 diode
R49342 N49341 N49342 10
D49342 N49342 0 diode
R49343 N49342 N49343 10
D49343 N49343 0 diode
R49344 N49343 N49344 10
D49344 N49344 0 diode
R49345 N49344 N49345 10
D49345 N49345 0 diode
R49346 N49345 N49346 10
D49346 N49346 0 diode
R49347 N49346 N49347 10
D49347 N49347 0 diode
R49348 N49347 N49348 10
D49348 N49348 0 diode
R49349 N49348 N49349 10
D49349 N49349 0 diode
R49350 N49349 N49350 10
D49350 N49350 0 diode
R49351 N49350 N49351 10
D49351 N49351 0 diode
R49352 N49351 N49352 10
D49352 N49352 0 diode
R49353 N49352 N49353 10
D49353 N49353 0 diode
R49354 N49353 N49354 10
D49354 N49354 0 diode
R49355 N49354 N49355 10
D49355 N49355 0 diode
R49356 N49355 N49356 10
D49356 N49356 0 diode
R49357 N49356 N49357 10
D49357 N49357 0 diode
R49358 N49357 N49358 10
D49358 N49358 0 diode
R49359 N49358 N49359 10
D49359 N49359 0 diode
R49360 N49359 N49360 10
D49360 N49360 0 diode
R49361 N49360 N49361 10
D49361 N49361 0 diode
R49362 N49361 N49362 10
D49362 N49362 0 diode
R49363 N49362 N49363 10
D49363 N49363 0 diode
R49364 N49363 N49364 10
D49364 N49364 0 diode
R49365 N49364 N49365 10
D49365 N49365 0 diode
R49366 N49365 N49366 10
D49366 N49366 0 diode
R49367 N49366 N49367 10
D49367 N49367 0 diode
R49368 N49367 N49368 10
D49368 N49368 0 diode
R49369 N49368 N49369 10
D49369 N49369 0 diode
R49370 N49369 N49370 10
D49370 N49370 0 diode
R49371 N49370 N49371 10
D49371 N49371 0 diode
R49372 N49371 N49372 10
D49372 N49372 0 diode
R49373 N49372 N49373 10
D49373 N49373 0 diode
R49374 N49373 N49374 10
D49374 N49374 0 diode
R49375 N49374 N49375 10
D49375 N49375 0 diode
R49376 N49375 N49376 10
D49376 N49376 0 diode
R49377 N49376 N49377 10
D49377 N49377 0 diode
R49378 N49377 N49378 10
D49378 N49378 0 diode
R49379 N49378 N49379 10
D49379 N49379 0 diode
R49380 N49379 N49380 10
D49380 N49380 0 diode
R49381 N49380 N49381 10
D49381 N49381 0 diode
R49382 N49381 N49382 10
D49382 N49382 0 diode
R49383 N49382 N49383 10
D49383 N49383 0 diode
R49384 N49383 N49384 10
D49384 N49384 0 diode
R49385 N49384 N49385 10
D49385 N49385 0 diode
R49386 N49385 N49386 10
D49386 N49386 0 diode
R49387 N49386 N49387 10
D49387 N49387 0 diode
R49388 N49387 N49388 10
D49388 N49388 0 diode
R49389 N49388 N49389 10
D49389 N49389 0 diode
R49390 N49389 N49390 10
D49390 N49390 0 diode
R49391 N49390 N49391 10
D49391 N49391 0 diode
R49392 N49391 N49392 10
D49392 N49392 0 diode
R49393 N49392 N49393 10
D49393 N49393 0 diode
R49394 N49393 N49394 10
D49394 N49394 0 diode
R49395 N49394 N49395 10
D49395 N49395 0 diode
R49396 N49395 N49396 10
D49396 N49396 0 diode
R49397 N49396 N49397 10
D49397 N49397 0 diode
R49398 N49397 N49398 10
D49398 N49398 0 diode
R49399 N49398 N49399 10
D49399 N49399 0 diode
R49400 N49399 N49400 10
D49400 N49400 0 diode
R49401 N49400 N49401 10
D49401 N49401 0 diode
R49402 N49401 N49402 10
D49402 N49402 0 diode
R49403 N49402 N49403 10
D49403 N49403 0 diode
R49404 N49403 N49404 10
D49404 N49404 0 diode
R49405 N49404 N49405 10
D49405 N49405 0 diode
R49406 N49405 N49406 10
D49406 N49406 0 diode
R49407 N49406 N49407 10
D49407 N49407 0 diode
R49408 N49407 N49408 10
D49408 N49408 0 diode
R49409 N49408 N49409 10
D49409 N49409 0 diode
R49410 N49409 N49410 10
D49410 N49410 0 diode
R49411 N49410 N49411 10
D49411 N49411 0 diode
R49412 N49411 N49412 10
D49412 N49412 0 diode
R49413 N49412 N49413 10
D49413 N49413 0 diode
R49414 N49413 N49414 10
D49414 N49414 0 diode
R49415 N49414 N49415 10
D49415 N49415 0 diode
R49416 N49415 N49416 10
D49416 N49416 0 diode
R49417 N49416 N49417 10
D49417 N49417 0 diode
R49418 N49417 N49418 10
D49418 N49418 0 diode
R49419 N49418 N49419 10
D49419 N49419 0 diode
R49420 N49419 N49420 10
D49420 N49420 0 diode
R49421 N49420 N49421 10
D49421 N49421 0 diode
R49422 N49421 N49422 10
D49422 N49422 0 diode
R49423 N49422 N49423 10
D49423 N49423 0 diode
R49424 N49423 N49424 10
D49424 N49424 0 diode
R49425 N49424 N49425 10
D49425 N49425 0 diode
R49426 N49425 N49426 10
D49426 N49426 0 diode
R49427 N49426 N49427 10
D49427 N49427 0 diode
R49428 N49427 N49428 10
D49428 N49428 0 diode
R49429 N49428 N49429 10
D49429 N49429 0 diode
R49430 N49429 N49430 10
D49430 N49430 0 diode
R49431 N49430 N49431 10
D49431 N49431 0 diode
R49432 N49431 N49432 10
D49432 N49432 0 diode
R49433 N49432 N49433 10
D49433 N49433 0 diode
R49434 N49433 N49434 10
D49434 N49434 0 diode
R49435 N49434 N49435 10
D49435 N49435 0 diode
R49436 N49435 N49436 10
D49436 N49436 0 diode
R49437 N49436 N49437 10
D49437 N49437 0 diode
R49438 N49437 N49438 10
D49438 N49438 0 diode
R49439 N49438 N49439 10
D49439 N49439 0 diode
R49440 N49439 N49440 10
D49440 N49440 0 diode
R49441 N49440 N49441 10
D49441 N49441 0 diode
R49442 N49441 N49442 10
D49442 N49442 0 diode
R49443 N49442 N49443 10
D49443 N49443 0 diode
R49444 N49443 N49444 10
D49444 N49444 0 diode
R49445 N49444 N49445 10
D49445 N49445 0 diode
R49446 N49445 N49446 10
D49446 N49446 0 diode
R49447 N49446 N49447 10
D49447 N49447 0 diode
R49448 N49447 N49448 10
D49448 N49448 0 diode
R49449 N49448 N49449 10
D49449 N49449 0 diode
R49450 N49449 N49450 10
D49450 N49450 0 diode
R49451 N49450 N49451 10
D49451 N49451 0 diode
R49452 N49451 N49452 10
D49452 N49452 0 diode
R49453 N49452 N49453 10
D49453 N49453 0 diode
R49454 N49453 N49454 10
D49454 N49454 0 diode
R49455 N49454 N49455 10
D49455 N49455 0 diode
R49456 N49455 N49456 10
D49456 N49456 0 diode
R49457 N49456 N49457 10
D49457 N49457 0 diode
R49458 N49457 N49458 10
D49458 N49458 0 diode
R49459 N49458 N49459 10
D49459 N49459 0 diode
R49460 N49459 N49460 10
D49460 N49460 0 diode
R49461 N49460 N49461 10
D49461 N49461 0 diode
R49462 N49461 N49462 10
D49462 N49462 0 diode
R49463 N49462 N49463 10
D49463 N49463 0 diode
R49464 N49463 N49464 10
D49464 N49464 0 diode
R49465 N49464 N49465 10
D49465 N49465 0 diode
R49466 N49465 N49466 10
D49466 N49466 0 diode
R49467 N49466 N49467 10
D49467 N49467 0 diode
R49468 N49467 N49468 10
D49468 N49468 0 diode
R49469 N49468 N49469 10
D49469 N49469 0 diode
R49470 N49469 N49470 10
D49470 N49470 0 diode
R49471 N49470 N49471 10
D49471 N49471 0 diode
R49472 N49471 N49472 10
D49472 N49472 0 diode
R49473 N49472 N49473 10
D49473 N49473 0 diode
R49474 N49473 N49474 10
D49474 N49474 0 diode
R49475 N49474 N49475 10
D49475 N49475 0 diode
R49476 N49475 N49476 10
D49476 N49476 0 diode
R49477 N49476 N49477 10
D49477 N49477 0 diode
R49478 N49477 N49478 10
D49478 N49478 0 diode
R49479 N49478 N49479 10
D49479 N49479 0 diode
R49480 N49479 N49480 10
D49480 N49480 0 diode
R49481 N49480 N49481 10
D49481 N49481 0 diode
R49482 N49481 N49482 10
D49482 N49482 0 diode
R49483 N49482 N49483 10
D49483 N49483 0 diode
R49484 N49483 N49484 10
D49484 N49484 0 diode
R49485 N49484 N49485 10
D49485 N49485 0 diode
R49486 N49485 N49486 10
D49486 N49486 0 diode
R49487 N49486 N49487 10
D49487 N49487 0 diode
R49488 N49487 N49488 10
D49488 N49488 0 diode
R49489 N49488 N49489 10
D49489 N49489 0 diode
R49490 N49489 N49490 10
D49490 N49490 0 diode
R49491 N49490 N49491 10
D49491 N49491 0 diode
R49492 N49491 N49492 10
D49492 N49492 0 diode
R49493 N49492 N49493 10
D49493 N49493 0 diode
R49494 N49493 N49494 10
D49494 N49494 0 diode
R49495 N49494 N49495 10
D49495 N49495 0 diode
R49496 N49495 N49496 10
D49496 N49496 0 diode
R49497 N49496 N49497 10
D49497 N49497 0 diode
R49498 N49497 N49498 10
D49498 N49498 0 diode
R49499 N49498 N49499 10
D49499 N49499 0 diode
R49500 N49499 N49500 10
D49500 N49500 0 diode
R49501 N49500 N49501 10
D49501 N49501 0 diode
R49502 N49501 N49502 10
D49502 N49502 0 diode
R49503 N49502 N49503 10
D49503 N49503 0 diode
R49504 N49503 N49504 10
D49504 N49504 0 diode
R49505 N49504 N49505 10
D49505 N49505 0 diode
R49506 N49505 N49506 10
D49506 N49506 0 diode
R49507 N49506 N49507 10
D49507 N49507 0 diode
R49508 N49507 N49508 10
D49508 N49508 0 diode
R49509 N49508 N49509 10
D49509 N49509 0 diode
R49510 N49509 N49510 10
D49510 N49510 0 diode
R49511 N49510 N49511 10
D49511 N49511 0 diode
R49512 N49511 N49512 10
D49512 N49512 0 diode
R49513 N49512 N49513 10
D49513 N49513 0 diode
R49514 N49513 N49514 10
D49514 N49514 0 diode
R49515 N49514 N49515 10
D49515 N49515 0 diode
R49516 N49515 N49516 10
D49516 N49516 0 diode
R49517 N49516 N49517 10
D49517 N49517 0 diode
R49518 N49517 N49518 10
D49518 N49518 0 diode
R49519 N49518 N49519 10
D49519 N49519 0 diode
R49520 N49519 N49520 10
D49520 N49520 0 diode
R49521 N49520 N49521 10
D49521 N49521 0 diode
R49522 N49521 N49522 10
D49522 N49522 0 diode
R49523 N49522 N49523 10
D49523 N49523 0 diode
R49524 N49523 N49524 10
D49524 N49524 0 diode
R49525 N49524 N49525 10
D49525 N49525 0 diode
R49526 N49525 N49526 10
D49526 N49526 0 diode
R49527 N49526 N49527 10
D49527 N49527 0 diode
R49528 N49527 N49528 10
D49528 N49528 0 diode
R49529 N49528 N49529 10
D49529 N49529 0 diode
R49530 N49529 N49530 10
D49530 N49530 0 diode
R49531 N49530 N49531 10
D49531 N49531 0 diode
R49532 N49531 N49532 10
D49532 N49532 0 diode
R49533 N49532 N49533 10
D49533 N49533 0 diode
R49534 N49533 N49534 10
D49534 N49534 0 diode
R49535 N49534 N49535 10
D49535 N49535 0 diode
R49536 N49535 N49536 10
D49536 N49536 0 diode
R49537 N49536 N49537 10
D49537 N49537 0 diode
R49538 N49537 N49538 10
D49538 N49538 0 diode
R49539 N49538 N49539 10
D49539 N49539 0 diode
R49540 N49539 N49540 10
D49540 N49540 0 diode
R49541 N49540 N49541 10
D49541 N49541 0 diode
R49542 N49541 N49542 10
D49542 N49542 0 diode
R49543 N49542 N49543 10
D49543 N49543 0 diode
R49544 N49543 N49544 10
D49544 N49544 0 diode
R49545 N49544 N49545 10
D49545 N49545 0 diode
R49546 N49545 N49546 10
D49546 N49546 0 diode
R49547 N49546 N49547 10
D49547 N49547 0 diode
R49548 N49547 N49548 10
D49548 N49548 0 diode
R49549 N49548 N49549 10
D49549 N49549 0 diode
R49550 N49549 N49550 10
D49550 N49550 0 diode
R49551 N49550 N49551 10
D49551 N49551 0 diode
R49552 N49551 N49552 10
D49552 N49552 0 diode
R49553 N49552 N49553 10
D49553 N49553 0 diode
R49554 N49553 N49554 10
D49554 N49554 0 diode
R49555 N49554 N49555 10
D49555 N49555 0 diode
R49556 N49555 N49556 10
D49556 N49556 0 diode
R49557 N49556 N49557 10
D49557 N49557 0 diode
R49558 N49557 N49558 10
D49558 N49558 0 diode
R49559 N49558 N49559 10
D49559 N49559 0 diode
R49560 N49559 N49560 10
D49560 N49560 0 diode
R49561 N49560 N49561 10
D49561 N49561 0 diode
R49562 N49561 N49562 10
D49562 N49562 0 diode
R49563 N49562 N49563 10
D49563 N49563 0 diode
R49564 N49563 N49564 10
D49564 N49564 0 diode
R49565 N49564 N49565 10
D49565 N49565 0 diode
R49566 N49565 N49566 10
D49566 N49566 0 diode
R49567 N49566 N49567 10
D49567 N49567 0 diode
R49568 N49567 N49568 10
D49568 N49568 0 diode
R49569 N49568 N49569 10
D49569 N49569 0 diode
R49570 N49569 N49570 10
D49570 N49570 0 diode
R49571 N49570 N49571 10
D49571 N49571 0 diode
R49572 N49571 N49572 10
D49572 N49572 0 diode
R49573 N49572 N49573 10
D49573 N49573 0 diode
R49574 N49573 N49574 10
D49574 N49574 0 diode
R49575 N49574 N49575 10
D49575 N49575 0 diode
R49576 N49575 N49576 10
D49576 N49576 0 diode
R49577 N49576 N49577 10
D49577 N49577 0 diode
R49578 N49577 N49578 10
D49578 N49578 0 diode
R49579 N49578 N49579 10
D49579 N49579 0 diode
R49580 N49579 N49580 10
D49580 N49580 0 diode
R49581 N49580 N49581 10
D49581 N49581 0 diode
R49582 N49581 N49582 10
D49582 N49582 0 diode
R49583 N49582 N49583 10
D49583 N49583 0 diode
R49584 N49583 N49584 10
D49584 N49584 0 diode
R49585 N49584 N49585 10
D49585 N49585 0 diode
R49586 N49585 N49586 10
D49586 N49586 0 diode
R49587 N49586 N49587 10
D49587 N49587 0 diode
R49588 N49587 N49588 10
D49588 N49588 0 diode
R49589 N49588 N49589 10
D49589 N49589 0 diode
R49590 N49589 N49590 10
D49590 N49590 0 diode
R49591 N49590 N49591 10
D49591 N49591 0 diode
R49592 N49591 N49592 10
D49592 N49592 0 diode
R49593 N49592 N49593 10
D49593 N49593 0 diode
R49594 N49593 N49594 10
D49594 N49594 0 diode
R49595 N49594 N49595 10
D49595 N49595 0 diode
R49596 N49595 N49596 10
D49596 N49596 0 diode
R49597 N49596 N49597 10
D49597 N49597 0 diode
R49598 N49597 N49598 10
D49598 N49598 0 diode
R49599 N49598 N49599 10
D49599 N49599 0 diode
R49600 N49599 N49600 10
D49600 N49600 0 diode
R49601 N49600 N49601 10
D49601 N49601 0 diode
R49602 N49601 N49602 10
D49602 N49602 0 diode
R49603 N49602 N49603 10
D49603 N49603 0 diode
R49604 N49603 N49604 10
D49604 N49604 0 diode
R49605 N49604 N49605 10
D49605 N49605 0 diode
R49606 N49605 N49606 10
D49606 N49606 0 diode
R49607 N49606 N49607 10
D49607 N49607 0 diode
R49608 N49607 N49608 10
D49608 N49608 0 diode
R49609 N49608 N49609 10
D49609 N49609 0 diode
R49610 N49609 N49610 10
D49610 N49610 0 diode
R49611 N49610 N49611 10
D49611 N49611 0 diode
R49612 N49611 N49612 10
D49612 N49612 0 diode
R49613 N49612 N49613 10
D49613 N49613 0 diode
R49614 N49613 N49614 10
D49614 N49614 0 diode
R49615 N49614 N49615 10
D49615 N49615 0 diode
R49616 N49615 N49616 10
D49616 N49616 0 diode
R49617 N49616 N49617 10
D49617 N49617 0 diode
R49618 N49617 N49618 10
D49618 N49618 0 diode
R49619 N49618 N49619 10
D49619 N49619 0 diode
R49620 N49619 N49620 10
D49620 N49620 0 diode
R49621 N49620 N49621 10
D49621 N49621 0 diode
R49622 N49621 N49622 10
D49622 N49622 0 diode
R49623 N49622 N49623 10
D49623 N49623 0 diode
R49624 N49623 N49624 10
D49624 N49624 0 diode
R49625 N49624 N49625 10
D49625 N49625 0 diode
R49626 N49625 N49626 10
D49626 N49626 0 diode
R49627 N49626 N49627 10
D49627 N49627 0 diode
R49628 N49627 N49628 10
D49628 N49628 0 diode
R49629 N49628 N49629 10
D49629 N49629 0 diode
R49630 N49629 N49630 10
D49630 N49630 0 diode
R49631 N49630 N49631 10
D49631 N49631 0 diode
R49632 N49631 N49632 10
D49632 N49632 0 diode
R49633 N49632 N49633 10
D49633 N49633 0 diode
R49634 N49633 N49634 10
D49634 N49634 0 diode
R49635 N49634 N49635 10
D49635 N49635 0 diode
R49636 N49635 N49636 10
D49636 N49636 0 diode
R49637 N49636 N49637 10
D49637 N49637 0 diode
R49638 N49637 N49638 10
D49638 N49638 0 diode
R49639 N49638 N49639 10
D49639 N49639 0 diode
R49640 N49639 N49640 10
D49640 N49640 0 diode
R49641 N49640 N49641 10
D49641 N49641 0 diode
R49642 N49641 N49642 10
D49642 N49642 0 diode
R49643 N49642 N49643 10
D49643 N49643 0 diode
R49644 N49643 N49644 10
D49644 N49644 0 diode
R49645 N49644 N49645 10
D49645 N49645 0 diode
R49646 N49645 N49646 10
D49646 N49646 0 diode
R49647 N49646 N49647 10
D49647 N49647 0 diode
R49648 N49647 N49648 10
D49648 N49648 0 diode
R49649 N49648 N49649 10
D49649 N49649 0 diode
R49650 N49649 N49650 10
D49650 N49650 0 diode
R49651 N49650 N49651 10
D49651 N49651 0 diode
R49652 N49651 N49652 10
D49652 N49652 0 diode
R49653 N49652 N49653 10
D49653 N49653 0 diode
R49654 N49653 N49654 10
D49654 N49654 0 diode
R49655 N49654 N49655 10
D49655 N49655 0 diode
R49656 N49655 N49656 10
D49656 N49656 0 diode
R49657 N49656 N49657 10
D49657 N49657 0 diode
R49658 N49657 N49658 10
D49658 N49658 0 diode
R49659 N49658 N49659 10
D49659 N49659 0 diode
R49660 N49659 N49660 10
D49660 N49660 0 diode
R49661 N49660 N49661 10
D49661 N49661 0 diode
R49662 N49661 N49662 10
D49662 N49662 0 diode
R49663 N49662 N49663 10
D49663 N49663 0 diode
R49664 N49663 N49664 10
D49664 N49664 0 diode
R49665 N49664 N49665 10
D49665 N49665 0 diode
R49666 N49665 N49666 10
D49666 N49666 0 diode
R49667 N49666 N49667 10
D49667 N49667 0 diode
R49668 N49667 N49668 10
D49668 N49668 0 diode
R49669 N49668 N49669 10
D49669 N49669 0 diode
R49670 N49669 N49670 10
D49670 N49670 0 diode
R49671 N49670 N49671 10
D49671 N49671 0 diode
R49672 N49671 N49672 10
D49672 N49672 0 diode
R49673 N49672 N49673 10
D49673 N49673 0 diode
R49674 N49673 N49674 10
D49674 N49674 0 diode
R49675 N49674 N49675 10
D49675 N49675 0 diode
R49676 N49675 N49676 10
D49676 N49676 0 diode
R49677 N49676 N49677 10
D49677 N49677 0 diode
R49678 N49677 N49678 10
D49678 N49678 0 diode
R49679 N49678 N49679 10
D49679 N49679 0 diode
R49680 N49679 N49680 10
D49680 N49680 0 diode
R49681 N49680 N49681 10
D49681 N49681 0 diode
R49682 N49681 N49682 10
D49682 N49682 0 diode
R49683 N49682 N49683 10
D49683 N49683 0 diode
R49684 N49683 N49684 10
D49684 N49684 0 diode
R49685 N49684 N49685 10
D49685 N49685 0 diode
R49686 N49685 N49686 10
D49686 N49686 0 diode
R49687 N49686 N49687 10
D49687 N49687 0 diode
R49688 N49687 N49688 10
D49688 N49688 0 diode
R49689 N49688 N49689 10
D49689 N49689 0 diode
R49690 N49689 N49690 10
D49690 N49690 0 diode
R49691 N49690 N49691 10
D49691 N49691 0 diode
R49692 N49691 N49692 10
D49692 N49692 0 diode
R49693 N49692 N49693 10
D49693 N49693 0 diode
R49694 N49693 N49694 10
D49694 N49694 0 diode
R49695 N49694 N49695 10
D49695 N49695 0 diode
R49696 N49695 N49696 10
D49696 N49696 0 diode
R49697 N49696 N49697 10
D49697 N49697 0 diode
R49698 N49697 N49698 10
D49698 N49698 0 diode
R49699 N49698 N49699 10
D49699 N49699 0 diode
R49700 N49699 N49700 10
D49700 N49700 0 diode
R49701 N49700 N49701 10
D49701 N49701 0 diode
R49702 N49701 N49702 10
D49702 N49702 0 diode
R49703 N49702 N49703 10
D49703 N49703 0 diode
R49704 N49703 N49704 10
D49704 N49704 0 diode
R49705 N49704 N49705 10
D49705 N49705 0 diode
R49706 N49705 N49706 10
D49706 N49706 0 diode
R49707 N49706 N49707 10
D49707 N49707 0 diode
R49708 N49707 N49708 10
D49708 N49708 0 diode
R49709 N49708 N49709 10
D49709 N49709 0 diode
R49710 N49709 N49710 10
D49710 N49710 0 diode
R49711 N49710 N49711 10
D49711 N49711 0 diode
R49712 N49711 N49712 10
D49712 N49712 0 diode
R49713 N49712 N49713 10
D49713 N49713 0 diode
R49714 N49713 N49714 10
D49714 N49714 0 diode
R49715 N49714 N49715 10
D49715 N49715 0 diode
R49716 N49715 N49716 10
D49716 N49716 0 diode
R49717 N49716 N49717 10
D49717 N49717 0 diode
R49718 N49717 N49718 10
D49718 N49718 0 diode
R49719 N49718 N49719 10
D49719 N49719 0 diode
R49720 N49719 N49720 10
D49720 N49720 0 diode
R49721 N49720 N49721 10
D49721 N49721 0 diode
R49722 N49721 N49722 10
D49722 N49722 0 diode
R49723 N49722 N49723 10
D49723 N49723 0 diode
R49724 N49723 N49724 10
D49724 N49724 0 diode
R49725 N49724 N49725 10
D49725 N49725 0 diode
R49726 N49725 N49726 10
D49726 N49726 0 diode
R49727 N49726 N49727 10
D49727 N49727 0 diode
R49728 N49727 N49728 10
D49728 N49728 0 diode
R49729 N49728 N49729 10
D49729 N49729 0 diode
R49730 N49729 N49730 10
D49730 N49730 0 diode
R49731 N49730 N49731 10
D49731 N49731 0 diode
R49732 N49731 N49732 10
D49732 N49732 0 diode
R49733 N49732 N49733 10
D49733 N49733 0 diode
R49734 N49733 N49734 10
D49734 N49734 0 diode
R49735 N49734 N49735 10
D49735 N49735 0 diode
R49736 N49735 N49736 10
D49736 N49736 0 diode
R49737 N49736 N49737 10
D49737 N49737 0 diode
R49738 N49737 N49738 10
D49738 N49738 0 diode
R49739 N49738 N49739 10
D49739 N49739 0 diode
R49740 N49739 N49740 10
D49740 N49740 0 diode
R49741 N49740 N49741 10
D49741 N49741 0 diode
R49742 N49741 N49742 10
D49742 N49742 0 diode
R49743 N49742 N49743 10
D49743 N49743 0 diode
R49744 N49743 N49744 10
D49744 N49744 0 diode
R49745 N49744 N49745 10
D49745 N49745 0 diode
R49746 N49745 N49746 10
D49746 N49746 0 diode
R49747 N49746 N49747 10
D49747 N49747 0 diode
R49748 N49747 N49748 10
D49748 N49748 0 diode
R49749 N49748 N49749 10
D49749 N49749 0 diode
R49750 N49749 N49750 10
D49750 N49750 0 diode
R49751 N49750 N49751 10
D49751 N49751 0 diode
R49752 N49751 N49752 10
D49752 N49752 0 diode
R49753 N49752 N49753 10
D49753 N49753 0 diode
R49754 N49753 N49754 10
D49754 N49754 0 diode
R49755 N49754 N49755 10
D49755 N49755 0 diode
R49756 N49755 N49756 10
D49756 N49756 0 diode
R49757 N49756 N49757 10
D49757 N49757 0 diode
R49758 N49757 N49758 10
D49758 N49758 0 diode
R49759 N49758 N49759 10
D49759 N49759 0 diode
R49760 N49759 N49760 10
D49760 N49760 0 diode
R49761 N49760 N49761 10
D49761 N49761 0 diode
R49762 N49761 N49762 10
D49762 N49762 0 diode
R49763 N49762 N49763 10
D49763 N49763 0 diode
R49764 N49763 N49764 10
D49764 N49764 0 diode
R49765 N49764 N49765 10
D49765 N49765 0 diode
R49766 N49765 N49766 10
D49766 N49766 0 diode
R49767 N49766 N49767 10
D49767 N49767 0 diode
R49768 N49767 N49768 10
D49768 N49768 0 diode
R49769 N49768 N49769 10
D49769 N49769 0 diode
R49770 N49769 N49770 10
D49770 N49770 0 diode
R49771 N49770 N49771 10
D49771 N49771 0 diode
R49772 N49771 N49772 10
D49772 N49772 0 diode
R49773 N49772 N49773 10
D49773 N49773 0 diode
R49774 N49773 N49774 10
D49774 N49774 0 diode
R49775 N49774 N49775 10
D49775 N49775 0 diode
R49776 N49775 N49776 10
D49776 N49776 0 diode
R49777 N49776 N49777 10
D49777 N49777 0 diode
R49778 N49777 N49778 10
D49778 N49778 0 diode
R49779 N49778 N49779 10
D49779 N49779 0 diode
R49780 N49779 N49780 10
D49780 N49780 0 diode
R49781 N49780 N49781 10
D49781 N49781 0 diode
R49782 N49781 N49782 10
D49782 N49782 0 diode
R49783 N49782 N49783 10
D49783 N49783 0 diode
R49784 N49783 N49784 10
D49784 N49784 0 diode
R49785 N49784 N49785 10
D49785 N49785 0 diode
R49786 N49785 N49786 10
D49786 N49786 0 diode
R49787 N49786 N49787 10
D49787 N49787 0 diode
R49788 N49787 N49788 10
D49788 N49788 0 diode
R49789 N49788 N49789 10
D49789 N49789 0 diode
R49790 N49789 N49790 10
D49790 N49790 0 diode
R49791 N49790 N49791 10
D49791 N49791 0 diode
R49792 N49791 N49792 10
D49792 N49792 0 diode
R49793 N49792 N49793 10
D49793 N49793 0 diode
R49794 N49793 N49794 10
D49794 N49794 0 diode
R49795 N49794 N49795 10
D49795 N49795 0 diode
R49796 N49795 N49796 10
D49796 N49796 0 diode
R49797 N49796 N49797 10
D49797 N49797 0 diode
R49798 N49797 N49798 10
D49798 N49798 0 diode
R49799 N49798 N49799 10
D49799 N49799 0 diode
R49800 N49799 N49800 10
D49800 N49800 0 diode
R49801 N49800 N49801 10
D49801 N49801 0 diode
R49802 N49801 N49802 10
D49802 N49802 0 diode
R49803 N49802 N49803 10
D49803 N49803 0 diode
R49804 N49803 N49804 10
D49804 N49804 0 diode
R49805 N49804 N49805 10
D49805 N49805 0 diode
R49806 N49805 N49806 10
D49806 N49806 0 diode
R49807 N49806 N49807 10
D49807 N49807 0 diode
R49808 N49807 N49808 10
D49808 N49808 0 diode
R49809 N49808 N49809 10
D49809 N49809 0 diode
R49810 N49809 N49810 10
D49810 N49810 0 diode
R49811 N49810 N49811 10
D49811 N49811 0 diode
R49812 N49811 N49812 10
D49812 N49812 0 diode
R49813 N49812 N49813 10
D49813 N49813 0 diode
R49814 N49813 N49814 10
D49814 N49814 0 diode
R49815 N49814 N49815 10
D49815 N49815 0 diode
R49816 N49815 N49816 10
D49816 N49816 0 diode
R49817 N49816 N49817 10
D49817 N49817 0 diode
R49818 N49817 N49818 10
D49818 N49818 0 diode
R49819 N49818 N49819 10
D49819 N49819 0 diode
R49820 N49819 N49820 10
D49820 N49820 0 diode
R49821 N49820 N49821 10
D49821 N49821 0 diode
R49822 N49821 N49822 10
D49822 N49822 0 diode
R49823 N49822 N49823 10
D49823 N49823 0 diode
R49824 N49823 N49824 10
D49824 N49824 0 diode
R49825 N49824 N49825 10
D49825 N49825 0 diode
R49826 N49825 N49826 10
D49826 N49826 0 diode
R49827 N49826 N49827 10
D49827 N49827 0 diode
R49828 N49827 N49828 10
D49828 N49828 0 diode
R49829 N49828 N49829 10
D49829 N49829 0 diode
R49830 N49829 N49830 10
D49830 N49830 0 diode
R49831 N49830 N49831 10
D49831 N49831 0 diode
R49832 N49831 N49832 10
D49832 N49832 0 diode
R49833 N49832 N49833 10
D49833 N49833 0 diode
R49834 N49833 N49834 10
D49834 N49834 0 diode
R49835 N49834 N49835 10
D49835 N49835 0 diode
R49836 N49835 N49836 10
D49836 N49836 0 diode
R49837 N49836 N49837 10
D49837 N49837 0 diode
R49838 N49837 N49838 10
D49838 N49838 0 diode
R49839 N49838 N49839 10
D49839 N49839 0 diode
R49840 N49839 N49840 10
D49840 N49840 0 diode
R49841 N49840 N49841 10
D49841 N49841 0 diode
R49842 N49841 N49842 10
D49842 N49842 0 diode
R49843 N49842 N49843 10
D49843 N49843 0 diode
R49844 N49843 N49844 10
D49844 N49844 0 diode
R49845 N49844 N49845 10
D49845 N49845 0 diode
R49846 N49845 N49846 10
D49846 N49846 0 diode
R49847 N49846 N49847 10
D49847 N49847 0 diode
R49848 N49847 N49848 10
D49848 N49848 0 diode
R49849 N49848 N49849 10
D49849 N49849 0 diode
R49850 N49849 N49850 10
D49850 N49850 0 diode
R49851 N49850 N49851 10
D49851 N49851 0 diode
R49852 N49851 N49852 10
D49852 N49852 0 diode
R49853 N49852 N49853 10
D49853 N49853 0 diode
R49854 N49853 N49854 10
D49854 N49854 0 diode
R49855 N49854 N49855 10
D49855 N49855 0 diode
R49856 N49855 N49856 10
D49856 N49856 0 diode
R49857 N49856 N49857 10
D49857 N49857 0 diode
R49858 N49857 N49858 10
D49858 N49858 0 diode
R49859 N49858 N49859 10
D49859 N49859 0 diode
R49860 N49859 N49860 10
D49860 N49860 0 diode
R49861 N49860 N49861 10
D49861 N49861 0 diode
R49862 N49861 N49862 10
D49862 N49862 0 diode
R49863 N49862 N49863 10
D49863 N49863 0 diode
R49864 N49863 N49864 10
D49864 N49864 0 diode
R49865 N49864 N49865 10
D49865 N49865 0 diode
R49866 N49865 N49866 10
D49866 N49866 0 diode
R49867 N49866 N49867 10
D49867 N49867 0 diode
R49868 N49867 N49868 10
D49868 N49868 0 diode
R49869 N49868 N49869 10
D49869 N49869 0 diode
R49870 N49869 N49870 10
D49870 N49870 0 diode
R49871 N49870 N49871 10
D49871 N49871 0 diode
R49872 N49871 N49872 10
D49872 N49872 0 diode
R49873 N49872 N49873 10
D49873 N49873 0 diode
R49874 N49873 N49874 10
D49874 N49874 0 diode
R49875 N49874 N49875 10
D49875 N49875 0 diode
R49876 N49875 N49876 10
D49876 N49876 0 diode
R49877 N49876 N49877 10
D49877 N49877 0 diode
R49878 N49877 N49878 10
D49878 N49878 0 diode
R49879 N49878 N49879 10
D49879 N49879 0 diode
R49880 N49879 N49880 10
D49880 N49880 0 diode
R49881 N49880 N49881 10
D49881 N49881 0 diode
R49882 N49881 N49882 10
D49882 N49882 0 diode
R49883 N49882 N49883 10
D49883 N49883 0 diode
R49884 N49883 N49884 10
D49884 N49884 0 diode
R49885 N49884 N49885 10
D49885 N49885 0 diode
R49886 N49885 N49886 10
D49886 N49886 0 diode
R49887 N49886 N49887 10
D49887 N49887 0 diode
R49888 N49887 N49888 10
D49888 N49888 0 diode
R49889 N49888 N49889 10
D49889 N49889 0 diode
R49890 N49889 N49890 10
D49890 N49890 0 diode
R49891 N49890 N49891 10
D49891 N49891 0 diode
R49892 N49891 N49892 10
D49892 N49892 0 diode
R49893 N49892 N49893 10
D49893 N49893 0 diode
R49894 N49893 N49894 10
D49894 N49894 0 diode
R49895 N49894 N49895 10
D49895 N49895 0 diode
R49896 N49895 N49896 10
D49896 N49896 0 diode
R49897 N49896 N49897 10
D49897 N49897 0 diode
R49898 N49897 N49898 10
D49898 N49898 0 diode
R49899 N49898 N49899 10
D49899 N49899 0 diode
R49900 N49899 N49900 10
D49900 N49900 0 diode
R49901 N49900 N49901 10
D49901 N49901 0 diode
R49902 N49901 N49902 10
D49902 N49902 0 diode
R49903 N49902 N49903 10
D49903 N49903 0 diode
R49904 N49903 N49904 10
D49904 N49904 0 diode
R49905 N49904 N49905 10
D49905 N49905 0 diode
R49906 N49905 N49906 10
D49906 N49906 0 diode
R49907 N49906 N49907 10
D49907 N49907 0 diode
R49908 N49907 N49908 10
D49908 N49908 0 diode
R49909 N49908 N49909 10
D49909 N49909 0 diode
R49910 N49909 N49910 10
D49910 N49910 0 diode
R49911 N49910 N49911 10
D49911 N49911 0 diode
R49912 N49911 N49912 10
D49912 N49912 0 diode
R49913 N49912 N49913 10
D49913 N49913 0 diode
R49914 N49913 N49914 10
D49914 N49914 0 diode
R49915 N49914 N49915 10
D49915 N49915 0 diode
R49916 N49915 N49916 10
D49916 N49916 0 diode
R49917 N49916 N49917 10
D49917 N49917 0 diode
R49918 N49917 N49918 10
D49918 N49918 0 diode
R49919 N49918 N49919 10
D49919 N49919 0 diode
R49920 N49919 N49920 10
D49920 N49920 0 diode
R49921 N49920 N49921 10
D49921 N49921 0 diode
R49922 N49921 N49922 10
D49922 N49922 0 diode
R49923 N49922 N49923 10
D49923 N49923 0 diode
R49924 N49923 N49924 10
D49924 N49924 0 diode
R49925 N49924 N49925 10
D49925 N49925 0 diode
R49926 N49925 N49926 10
D49926 N49926 0 diode
R49927 N49926 N49927 10
D49927 N49927 0 diode
R49928 N49927 N49928 10
D49928 N49928 0 diode
R49929 N49928 N49929 10
D49929 N49929 0 diode
R49930 N49929 N49930 10
D49930 N49930 0 diode
R49931 N49930 N49931 10
D49931 N49931 0 diode
R49932 N49931 N49932 10
D49932 N49932 0 diode
R49933 N49932 N49933 10
D49933 N49933 0 diode
R49934 N49933 N49934 10
D49934 N49934 0 diode
R49935 N49934 N49935 10
D49935 N49935 0 diode
R49936 N49935 N49936 10
D49936 N49936 0 diode
R49937 N49936 N49937 10
D49937 N49937 0 diode
R49938 N49937 N49938 10
D49938 N49938 0 diode
R49939 N49938 N49939 10
D49939 N49939 0 diode
R49940 N49939 N49940 10
D49940 N49940 0 diode
R49941 N49940 N49941 10
D49941 N49941 0 diode
R49942 N49941 N49942 10
D49942 N49942 0 diode
R49943 N49942 N49943 10
D49943 N49943 0 diode
R49944 N49943 N49944 10
D49944 N49944 0 diode
R49945 N49944 N49945 10
D49945 N49945 0 diode
R49946 N49945 N49946 10
D49946 N49946 0 diode
R49947 N49946 N49947 10
D49947 N49947 0 diode
R49948 N49947 N49948 10
D49948 N49948 0 diode
R49949 N49948 N49949 10
D49949 N49949 0 diode
R49950 N49949 N49950 10
D49950 N49950 0 diode
R49951 N49950 N49951 10
D49951 N49951 0 diode
R49952 N49951 N49952 10
D49952 N49952 0 diode
R49953 N49952 N49953 10
D49953 N49953 0 diode
R49954 N49953 N49954 10
D49954 N49954 0 diode
R49955 N49954 N49955 10
D49955 N49955 0 diode
R49956 N49955 N49956 10
D49956 N49956 0 diode
R49957 N49956 N49957 10
D49957 N49957 0 diode
R49958 N49957 N49958 10
D49958 N49958 0 diode
R49959 N49958 N49959 10
D49959 N49959 0 diode
R49960 N49959 N49960 10
D49960 N49960 0 diode
R49961 N49960 N49961 10
D49961 N49961 0 diode
R49962 N49961 N49962 10
D49962 N49962 0 diode
R49963 N49962 N49963 10
D49963 N49963 0 diode
R49964 N49963 N49964 10
D49964 N49964 0 diode
R49965 N49964 N49965 10
D49965 N49965 0 diode
R49966 N49965 N49966 10
D49966 N49966 0 diode
R49967 N49966 N49967 10
D49967 N49967 0 diode
R49968 N49967 N49968 10
D49968 N49968 0 diode
R49969 N49968 N49969 10
D49969 N49969 0 diode
R49970 N49969 N49970 10
D49970 N49970 0 diode
R49971 N49970 N49971 10
D49971 N49971 0 diode
R49972 N49971 N49972 10
D49972 N49972 0 diode
R49973 N49972 N49973 10
D49973 N49973 0 diode
R49974 N49973 N49974 10
D49974 N49974 0 diode
R49975 N49974 N49975 10
D49975 N49975 0 diode
R49976 N49975 N49976 10
D49976 N49976 0 diode
R49977 N49976 N49977 10
D49977 N49977 0 diode
R49978 N49977 N49978 10
D49978 N49978 0 diode
R49979 N49978 N49979 10
D49979 N49979 0 diode
R49980 N49979 N49980 10
D49980 N49980 0 diode
R49981 N49980 N49981 10
D49981 N49981 0 diode
R49982 N49981 N49982 10
D49982 N49982 0 diode
R49983 N49982 N49983 10
D49983 N49983 0 diode
R49984 N49983 N49984 10
D49984 N49984 0 diode
R49985 N49984 N49985 10
D49985 N49985 0 diode
R49986 N49985 N49986 10
D49986 N49986 0 diode
R49987 N49986 N49987 10
D49987 N49987 0 diode
R49988 N49987 N49988 10
D49988 N49988 0 diode
R49989 N49988 N49989 10
D49989 N49989 0 diode
R49990 N49989 N49990 10
D49990 N49990 0 diode
R49991 N49990 N49991 10
D49991 N49991 0 diode
R49992 N49991 N49992 10
D49992 N49992 0 diode
R49993 N49992 N49993 10
D49993 N49993 0 diode
R49994 N49993 N49994 10
D49994 N49994 0 diode
R49995 N49994 N49995 10
D49995 N49995 0 diode
R49996 N49995 N49996 10
D49996 N49996 0 diode
R49997 N49996 N49997 10
D49997 N49997 0 diode
R49998 N49997 N49998 10
D49998 N49998 0 diode
R49999 N49998 N49999 10
D49999 N49999 0 diode
R50000 N49999 N50000 10
D50000 N50000 0 diode
.op
.control                                    ; begin of control section
<<<<<<< HEAD
run                                         ; run the .tran command
=======
run                                         ; run the .op command
print N0
>>>>>>> 94f60a3 (update)
print N50000
.endc 
.end