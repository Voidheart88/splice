Vin 1 0 10
R1 1 2 1000
E1 3 0 1 0 1.0
.op
.end